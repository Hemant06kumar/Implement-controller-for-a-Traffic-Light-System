%PDF-1.7
%����
9 0 obj
<<
/Ordering (Identity)
/Registry (Adobe)
/Supplement 0
>>
endobj
11 0 obj
<<
/Filter /FlateDecode
/Length 17
>>
stream
H�:�$� ��` � �
endstream
endobj
12 0 obj
<<
/Filter /FlateDecode
/Length 933
/Subtype /CIDFontType0C
>>
stream
H�|�mLSW������r����=검�4$��� '#��0-�.`os{�F�hXa8�"-���$��:ƲQ�f~ �^>,qƹ}Y���#��vo�%K��|��������OIl�D�$�܁�:�s_~��Do�$�{�U^��1(g�b��$�ތX�ƫ8���hoP/��mhg�R�l8�<B��:�H�IRdN�[l�kܼW�*��'	�2(,-��Z�V{Z��Z�֒`��li��������/������.J>Qrɼ{7���ik?�x?/���~���N^.��!(�%�d��揹�n ����F�/��Tr�J�\^�Uq�S��^�,	��u����ǃ��=��VY�����%�"⟥WtD7q�l"�61�#I�k�T4/�A��>�O�Q�G%OY�㳸��"]�:��J)�`��JH%��BF#���k�'�^�1K��Z(�`dm{��$��Yd�/ӵ�'O�0�L)Hi������=+uo���A�L�v��B��r��k�����VGcCK������������
���t<�0�� �0�#|B�нȷ?���Mt�g�=��
Ǻt��e�I_�d��q�i����l��6{ei��K�R���q���DG��	��b�RR(,�x�8����L�/�Z-����7ߋ}�C���W�,t��G5�c0Q�������ڕ[&.q�C�C�nn�ꢯ3X�9x>�m�������i.:nu|�`��'У8yj�n� +:I�	|67�I��o0��[���������w7�v�9m��|�.+�u�_�m�~��!03;4�@��!$����+_�t�|;����Wkc�Q����v��8��Au�S�5>�	���	��(��O@Kd"z%l���6���#T��5����l�J�%� W?��
endstream
endobj
10 0 obj
<<
/Ascent 1008
/CIDSet 11 0 R
/CapHeight 651
/Descent -360
/Flags 6
/FontBBox [-317 -360 1684 1008]
/FontFamily (Minion Pro Cond)
/FontFile3 12 0 R
/FontName /KTNQSD+MinionPro-BoldCn
/FontStretch /Condensed
/FontWeight 700
/ItalicAngle 0
/StemV 124
/Type /FontDescriptor
/XHeight 442
>>
endobj
8 0 obj
<<
/BaseFont /KTNQSD+MinionPro-BoldCn
/CIDSystemInfo 9 0 R
/DW 1000
/FontDescriptor 10 0 R
/Subtype /CIDFontType0
/Type /Font
/W [0 [500 195 267 346] 4 5 466 6 [730 667 226] 9 10 328 11 [385 577 248 309 248 303] 17 26 466 27 28 248 29 [554 577 554 383 719 633 588 583 668 532 510 631 697 346 332 634 504 801 656 654 554 651 610 471 561 655 638 879 617 595 553 325 305 325 559 500 226 439 500 394 510 415 305 454 514 275 271 486 261 782 527 488 506 502 379 364 318 512 437 642 454 439 415 327 245 327 577 267] 97 98 466 99 [168] 100 101 466 102 [464 466 179 418 449] 107 108 276 109 110 542 111 [504 480 473 248 477 384 236 440 418 449 899 1041 383] 124 136 400 137 [908 812 322 516 655 893 344 640 276 287 493 716 532 324 577 504 465 676 730 577 552 728 577 245 323 502 730 324 312 577 486 577 324 696] 171 176 633 177 [585] 178 181 532 182 185 346 186 [656] 187 191 654 192 [471] 193 196 655 197 198 595 199 [553] 200 205 439 206 [395] 207 210 415 211 214 276 215 [527] 216 220 488 221 [364] 222 225 512 226 227 439 228 [415 506 500 466 418] 233 238 730 239 [633 930 628 600 676 656 697 560 480 601 593 500 966 711 445 276 511 520 516 519 527 321 376 683 1012 889 861 719 791 570 1059 1064 809 800 1036 808 861 798 542 537 775 542 595 548 845 676 785 795 540 764] 289 290 540 291 [587 806 807] 294 298 466 299 [842 439 764 563 536 513 577 481 458 553 606 319 312 554 458 686 554 569 503 570 545 427 504 556 554 725 548 511 484] 328 329 606 330 [319 572 504 552 606 515 434 854 722 776 275 606 631 632] 344 345 255 346 347 381 348 [516 351 440 412 466 388 494 422 470 491 479 466 550 486 494 497 520 493 494 498 701 1014 697 496 351 461 455 485 453 497 462 486 493 496 476 460 566 475 502 466 563 481 503 464] 392 411 490 412 [322 362 368] 415 416 301 417 [321 382 209 208 558 384 344 275 278 235] 427 436 324 437 438 187 439 440 324 441 [259] 442 443 237 444 453 324 454 455 187 456 457 324 458 [259] 459 460 237 461 470 324 471 472 187 473 474 324 475 [259] 476 477 237 478 487 324 488 489 187 490 491 324 492 [259] 493 494 237 495 497 606 498 [454 469 407 554] 502 507 633 508 [1058 813] 510 512 633 513 520 697 521 [566 697] 523 526 687 527 [640 687 598 681] 531 532 652 533 534 877 535 536 631 537 540 687 541 542 504 543 [271] 544 545 846 546 [719 908 504 267] 550 551 449 552 553 276 554 [309 383] 556 557 327 558 559 325 560 561 328 562 [248] 563 564 570 565 [595 571 730 511 389 489 681 554 516 596 687 510 532] 578 580 633 581 [664] 582 585 583 586 [668] 587 590 532 591 [531] 592 596 631 597 [697] 598 602 346 603 [332 634] 605 608 504 609 [801] 610 613 656 614 616 654 617 [655] 618 620 610 621 [471 473] 623 624 471 625 626 561 627 632 655 633 636 879 637 639 595 640 641 553 642 [812] 643 644 1012 645 646 439 647 [440 490] 649 652 394 653 [510] 654 658 415 659 663 454 664 [514] 665 668 276 669 [274 486] 671 673 261 674 [311 782] 676 679 527 680 682 488 683 [493] 684 686 379 687 [364 367] 689 690 364 691 692 318 693 695 512 696 [515] 697 698 512 699 702 642 703 705 439 706 707 415 708 [640 400] 710 711 500 712 724 400 725 728 563 729 [722] 730 734 563 735 [582] 736 737 513 738 [515] 739 740 513 741 [577] 742 750 481 751 755 553 756 [606] 757 760 319 761 [471] 762 765 319 766 [312 554] 768 771 458 772 [479 686] 774 778 554 779 785 569 786 [572 569] 788 790 545 791 792 427 793 [426] 794 795 427 796 797 504 798 804 556 805 [557] 806 807 556 808 811 725 812 816 511 817 819 484 820 [400 401 400] 823 824 401 825 [407 401] 827 830 400 831 [401] 832 833 400 834 [633 588 496 596 532 553 697 651 346 634 636 801 656 576 654 679 554 555 561 603 723 617 714 687 633 532 697] 861 862 346 863 [654] 864 865 603 866 [687] 867 873 633 874 882 881 883 887 633 888 895 532 896 901 697 902 910 938 911 914 697 915 926 346 927 932 687 933 941 960 942 945 687 946 953 654 954 [554 346] 956 963 603 964 [346 332 823 898 706 621 588 694 633 578 588 490 614 532 892 496] 980 981 698 982 [621 606 801 697 654 681 554 583 561 504 501 468 476 393 363 495 482 264 477 473 504 452 392 488 487 489 430 452 572 448 567 611 384 487 471 562 623 395 489 669 525 447 504 393 495] 1027 1028 264 1029 [488] 1030 1031 452 1032 [611 264 452] 1035 1042 504 1043 1048 393 1049 1056 495 1057 1064 264 1065 1070 488 1071 1078 452 1079 1086 611 1087 1088 504 1089 1090 393 1091 1092 495 1093 1094 264 1095 1096 488 1097 1098 452 1099 1100 611 1101 1108 504 1109 1116 495 1117 1124 611 1125 1130 504 1131 1135 495 1136 1141 264 1142 1145 452 1146 1147 487 1148 [452] 1149 1153 611 1154 [504 452] 1156 1159 251 1160 1177 400 1178 1179 424 1180 [400 588 726 617 694 643 925 928 694 845 571 584 900 615 439 481 485 387 467 415 709 403] 1202 1203 537 1204 [496 473 600 534 488 532 506 394 424 439 670 454 540 501 759 760 554 696 465 420 710 498 415 491 387 420 364 275 276 271 648 703 517 496 445 531 668 544 646 488 615 449 451 365 422 309 432 865 974 1124 1133 957 457 603 623 830 1006 806 1408 1744 1095 643 566 821 836 906 1602 1675 1584 427 892] 1275 1276 745 1277 [465 619 734 427 346 566 892] 1284 1287 400 1288 [654 655 499 525] 1292 1293 466 1294 1305 633 1306 1313 532 1314 1315 346 1316 1327 654 1328 1334 655 1335 1337 595 1338 1349 439 1350 1357 415 1358 1359 276 1360 1366 488 1367 1371 499 1372 1373 512 1374 1378 525 1379 1381 439 1382 1393 601 1394 1401 593 1402 1413 563 1414 1421 481 1422 1423 319 1424 1436 569 1437 1444 556 1445 1447 511 1448 1457 400 1458 [372] 1459 1480 400 1481 [563 536 513 577 481 458 553 606 319 312 554 458 686 554 569 503 570 545 427 504 556 554 725 548 511 484] 1507 1508 606 1509 [572 504 552 606 515 434 722 776 631] 1518 1521 563 1522 [722] 1523 1528 563 1529 1530 513 1531 [515] 1532 1533 513 1534 [577] 1535 1543 481 1544 1548 553 1549 [606] 1550 1558 319 1559 [312 554] 1561 1564 458 1565 [479 686] 1567 1571 554 1572 1578 569 1579 [572 569] 1581 1583 545 1584 1585 427 1586 [426] 1587 1588 427 1589 1590 504 1591 1597 556 1598 [557] 1599 1600 556 1601 1604 725 1605 1609 511 1610 1612 484 1613 1624 563 1625 1632 481 1633 1634 319 1635 1647 569 1648 1655 556 1656 1658 511 1659 [473 367 561 318 309 195 400 168 248 319 168] 1670 1671 103 1672 [477 563 777 916 312 226 466 480 466 490 466 487 465 490]]
>>
endobj
7 0 obj
[8 0 R]
endobj
13 0 obj
<<
/Filter /FlateDecode
/Length 255
>>
stream
H�\��j�0��~
�Cqw;�@i7�aX�pl%3,�q�C�~�:����'����֚�=8�a��XpvKP=�Ʋ�mT܉~5I�xw�qj��X]�H�9��z<2�4cG8|]�#�n��'�
h�8�F/ҿ�	�����7q=%�_���*�2/����K�A�Y]�h�~N�0��_�1��A}�@�e�.��h��2݈JA$*�*�y�s&A$2=��wߦ�#�ݚZBH��dg3b,ޏ흇���` �}
endstream
endobj
6 0 obj
<<
/BaseFont /KTNQSD+MinionPro-BoldCn
/DescendantFonts 7 0 R
/Encoding /Identity-H
/Subtype /Type0
/ToUnicode 13 0 R
/Type /Font
>>
endobj
20 0 obj
<<
/Filter /FlateDecode
/Length 21
>>
stream
H�:� 
,���(  =�
endstream
endobj
21 0 obj
<<
/Filter /FlateDecode
/Length 2413
/Subtype /CIDFontType0C
>>
stream
H�|�kPS��O��=V�����s4'�u�����"2nU�Y��V�@��$$�$��K8	!B.r�1rQ��cWƶvUv�-������u[�N�c��9�Kg:�/��9�y�������p8�WS���%��&S�T���W{T
I��]�H�Ժ�!��C����1������WC���_P�?���Bm�ycݪc6 ь �Exȏ�κ�U�4E"U�d:c�Jm�ȊKt��		��e��p��[�5>\��+ڲiӦp��[Ea-Q�Q���iE)�B�F�҈uR�F�n�B�֊4R�TS�>|y�L+��t%R�H�,˘��D�ӈ%�2�F.R�+����Q"�R�h�r�2���1�"�R���
O)TU(u�T���l�Z*�.�H���[�'��� �#�ً �QHZ��A"�5Y��e�<�d"M�tp���u䟢����Fˣ�䊸~��`
���e��n���s�Tc܋���g j�����n�?���w����
��pG��v�L�㥴���r��H�����j��3F	�w�m�0DJ�m�mM�V �Z�B
K�����Nh��0>IMRF�}���|�r�R���sյξjB�m�'��)�9�w�#�ك�v�����+e��u�	gC`���� ��.��mU�DWUG�/��,eWR�3����������Fk]��2wN�C0SA��+��xF}Z�D�V�j�&L5�>�kr	�g�:�h���م��"
��r���=b�P�2~��<4
u�Z�������EPW[g7����s�ݣ=�)o��T�3�<���8Iq!�d�\�x�{�vid�X<N�{\�.�st�,q�g��|��T�-�29Dj~��$�����]�q�攐�ƨn��&9g ��H*���e�<%��?���Og:�px��'S�7��ye�RBVR����w߄��<�&�w�/c}9�F��D4ɚ%��s��8��)Ε�1(�љ7Z��_C��ꠀ?�*q�F�oݤ������:� ��ฅ�������y�׹���oZ�9O��������#Z�i��c�4�<�]��]��F��ܩ됴#K�����ǭ�(Ya�Wb���͟���彩[�a�U����<�9�*�-z�??O�Q���R�	�xʿ8�+WzN�[6��i����)Q�AQ�W�lr۫}�~�x��,�WQC�լǲo��Wa�#�������-,S5��BS�����Φv&��'_�=�U����A��{�Ջ��i�E0՟���P,k&
��K�Cg��~�s��PS���*��ٗ;}�����3����9���%�/B��s�9c�ERqA�����7<?�����
�^թ�\U��d[K�R �DrlL"� (r��b���܃�ĨfA��L�M�dx�z&�D�r�b����[p>�<�<#-V�I�A��+nA�H�m>�U-YVTf�Mi] >���Ȱ�;-�o�9��b�9���Q@vu2������tl%����0�e���K��q��Լ�Nf�Q��m�G�c��v��\�jM���2����Z�^A,��*z���9h9�RwҞ��
�f�g1\��u�d�h}��C�Ĉ� A��t[��}C/�� o���K8�u�3���cI[��������R6���=�"�dP��N����\h�T��f�8l:d>�R]�o���T���0U%C�$71�
��z=��]2;-���r�R�$��un�x$<I��^��N��;4�o����p\��:���
���Ac��%*Y��	|��k��[Z�{�X*�5��.2���,̣��; ݐn̬CU`���ض��1�<�^�� �Ǆ�D��}���!/��	|{����0�mu���D����3��\?J��׈�Oh���F�W�xu�o����z`�A��� ����:\�u�r1Z2H���wd���X������v��]�K�&=M~':�9=:��ӌ���L|PN���LP��9����y$�.��j�Z���� =����Ig�ļ��\�)*�Y�?��	��ɢ�d����Y�<�����_d�� �T������ ��hH�-�\v�,�h�����ʭ���~}�uro�����������-�}�� ?EhXph��h���2�hҖ������hv����R�&�
�X�N�<m����gyIr;sCG�o��������}m����_�[����+�z�}�|���z�z|qv|kwv��|l�n������������5��!�գġ��� 
�&�
~��N����������}�|��I����%��������	�F�_	��
��W�0 �֖X
endstream
endobj
22 0 obj
<<
/Filter /FlateDecode
/Length 317
>>
stream
H�\�ۊ�0�{�b.ۋ�*�Pz /���� ��]a�!��~c�҅(|$�df⟪s����w3��g�z%O����o��d/��_��|\/��C���+
�?��4��6G9����7#���F��S�%��k����*K��ٍ^��L��U����1+>�9���%O�luc��(���Qz���0GXۉ�Ƹ�]QP���Nq�O���)�����=�B	�A)t�2(��Kq^|�N�:CW���BrH�P�� �%8=�]�5Y�f{Kώ��1���.���?߈5٨��~ |Ԡ�
endstream
endobj
27 0 obj
<<
/Filter /FlateDecode
/Length 23264
/Length1 50536
/Type /Stream
>>
stream
x��\UU�7�.{�s� DT8�xE@��@@QDTLS��`܆��L��{�h��9���k��Լ����VcMW�Ɇ�e���~�����f���~��y>�s����k���~k�J�G�Grr֘�Wn\'�t*zۏHLJ^�^e9!K��~�����юKg	yt!o���0y�G	9>.�i������1~|nIN�忕��bB�S���WkL6B�\$����(�������9X� KO��6�xn�*��%B�+S_���gr���xޯ�Z��4��
K���Sp�6xfqYnζ�_'d���+əS���%�/G��4�$���.'����!�e�U��d��)��W�z�8�;j	1���bSj7>�f��;�{j&���=~t_Z�@գ恸5��3�� �?�t�G%&�E�x�"1��{F�d���N���r��#*zz��qb\�����c��f�f�1�盧�� ��bbzAR�#�S��S	�b��8?�_ ���,L�X�(�H2;�C'�]$���y�*) K�M���@k-ګ���^��I������Uq���+�YR��}2�����U$��'BF����M
�}d$�j����d>�,�!RG��I�9JVЙ��=I��SA�䯐�_�>�ǳU�M����0`�!�A?��!�Z	4�~��3A�**h~Tx�4��.8����q��xz�7A7�`���ِ�I��B`Y�XV�׳� 3��;��E��I2h:в8��z�����@��7�MH�s�@�v��h,#�Y��y]%%�T��ws�T�O��w+��.'Aq ��x�`�L��c3���,����è>�=���(����t�Tj�Az��@�k%5sȬFz,�E�?p�X@�{�d�t �ɸ����X�N��k�����5JH`;${�H�1f��sإ��.��筠�R��U��\@�I����9	b��VD�Nfb�!�=G�.���'_¬��k�kM���s��F�Bȳ�d?fχ�灃ش���ȫ�����)���{9Y�U��ԛ t&�����n���%��T�l$�E)�����"\�J.`�~��:��{.{;�'�!
n&&�ȗ�C�t-�=M�_�̀{id�G��ۀ���@7ڍu�CD�s��P��F3J�ӝ4�f�O��'Q̉ty���m��J� r�ð�x��at<y�F.�b��
[�9ZIOo���5�䠜��nB��ZƑ�er�Č�l�u41c�89b���T�3 |})l��H]�"Җ`�a$�^u���8C��˝o�~2�4lD��Yi�e,���x���jXQ5��,����I��V|g�7�X��:��Vف�t���@�02�L�>��r�F�
��I�p �S���<��O�4��o"z�Cx�pw�@�B2�UF�u��-<���	C��T(9�%�눑��W� ��;���p���
D,#���������5�6?D�uRR���b�h/ �܋qid���p�?	_: �$+���I9ʁт��1f�W_�$$*bC(�N~�"Dc�2Y��}g]��$5衯5�1��ϓō7؅oU��J����'^���c��l���C=������zĆ�ѷY�T\ǣġLC�4`�&�u�ף���F��ޣ��gt.ds��E��D�6�	��#��G���x���
_&�b�nX�ˈ��;�/\'`tW2�:�{���xy�{�2=@	}���1b��(I�,�+�����CSV��u΃Ѓ�'���!� �Q���Á0޸�xyׇ ;�����&y��j�\�\� �{�sd/5��ג����E� �!�����L��"R��v<���2�L �4�᤟V��տJ2@��C��י44��8�c���)����)�U�m�-�m��˻�r�S��yZ>݆�,Wk�=��R����'`�B�>��rX�0�z�=�HD�A����$ڎD!��QF���%A�?��^���4�@䝄��(��3�N"N�ӑ���h8�O!�mǳl��A�7�u��9�0�"b҇0+B��I\��:���dz~9�{��%�]��;�r���gfuc���@:+��py�Q�o�KA�%��e6gĬ��ٔ(Cd��l�N�@X�@�	��#b�("/h�g���Pr�q��
w��MDf�Y��"��,FFg����Z/֋��&�+ε2�p�s�saê�U���Fc>��瘆8�Άuz������{څ��*��l�)����}��
��.�O�+���~8����tbN����{�_��,�H�_ #�'1���^���+��[k7��\��A��B�w��&��d��o@��M(�~�^9
��~��'�Y���UP=	9�B���W��.���o�Q�8�yGù�6���Vfa�q�{���uvSc�^چ,r��ѝ�<�_�y��î��oȓ�Hjü��ATn/�@<z�3ܝ�'!�B$ꅑ�#pc��|�h�TW�ڈ����:�w�p_X1�� 2	+�~5l}����pv'����r���z[Om�Xj]� �h|&�h��\��Bܽ�^���)kc��u���O��<��'�DO��w� A�qߵ�*G�"2ʃ2'Jq�r�"���[�\�V�[@v���{$�=���.X���Lt�~�:���Y&4k�4�tی�.�p[Od���� ��)���A�Z�l/�ѫ���?:DNs������tߧ�\�n�"
� ޢ`d�T�]�"#H6��^F�e�lFù+�9�	�*�Ш�7��i�;��w�Y'�	5C���My��]��V?Ěd��ʾd�<#]ke���F%��4��dߣ؈���3/
���F�ru,��An?���EMψ�Ƙ;߻����
�t8��\��9�u�ܾX��~F���P�B��U~X�o�uJ���|"��� �v�	��k��\���;b�D��^]挀fχ���3�i����ϡ�C��<��AD�s�?��(�gf�ι�N{�� �wF���.���p����Ӆ�g��Èvr7�9���q@kx�>�R��"V�évp�-�t"b�p�k9��0o&��@>�Y8]� C,N�^��"Q�{�L�i�	���a=�q��S�hd�=��E��(D����F���T���V�b`�tJr��@�9t��W!à۞��Q�A�&�X���dq�} ��'qVY���m_m�F�$6%eJx��1��<�ъ_��NG�� "�ā� \���-hꄨ<Ҋ!=X;�&����wnBJND�(D�x�N��Z�L?��x��E��p2�$U��D\�D�O����3z?ҏ�E-�Q}��ػ��#�Y��xw�}a9�%������jڍv���GEf��*@�Z�]�ZF�tH[\��9yhD��;X�Z�v<�ϔ'�T�Μ~I���8yd�c8N���Y4�u�<��� |�?�3����������
h'\�����ͫ�s��U�d�3�4Q�չD��������㊄A���'���DTqߡĠ�G�xB��W ���A��=1?��֏ɷ���st~e��Ng'�I��j�O{^��4��#<��r	u~#�f���:����d��7��
~/n~��q$��)��T��D�?ȝ�����>)���7"��'��22�o'���0<p��~�3�0���|��� ����6D�	?�X>f
(}E�SQ�'\�2'���0��T�sW�N�-u�x(b�x��XY�ab�l2����9�-FuE����)X{,<~*���*bu:�_�"��v�gsw�����?�2�i\���F�����W|
����P�xW�2eJg�W��Z#�V�&��(�(�(Y(���$JJ���Q@)GIC� �}�^E��e2���(�)�O�[|h��94~Srw�6YP�Ѫ�a�"c&w����%��]���c�
���{C ,%{j{D�ؒ;qI�3����aw�T�<b\� R
��H��H"l2�	��¾*$�&s�{�yB��\'�������?^�{}���h�T�#ǎt�������q�f;�L��3�ŭ�nr�'����:j���l��:q��~?�0�W"�?���������m�]h��%�33Mq�n�'%�gb��j��L���-t����Ҟ?��Klm}`��j|{�3G��(4��h���?�S?ٶ�ڗlA�#���1B����H8�!�r����*�Y�(3��S�lkr�*ۊ�粇�7Q���z����[��_����7W�?�������'�7W󛋔�otV��ȿ�Snt��}�~w���[��u��X~-���ׁ�:���:/�9���__�S��ȯ��t��/۩������t~����??�?�4H���4��������[�������F��Z���k��Z�����K��4�_����X�wu���_��y����O}�=�S��6�7VE�o��u��]����5�����[��S:?��:E�ǁ�x ?f�G_>����G�W_>�_^�9����SG�C:i#�]�������\/���<~ ��ɇ�����|������:��?ߣ�gw������>��]~�3]�.?�_;{���������:Z�۷�������� �����ʷ��I,�ηx�͛���:��k�~�F����F�?�z�0b��a]���~�!NY�����q�?~����k!����1p�X _��W�cu_����+��
�/��2�?��O}T�K��#:_���ԇ3�b�/��>�@]���!�A�����t>[�t^]eS�}yu-%q��*�:�T���8�B��y���J3ղ�����Z��K��b�?�g�(���3����<O��C�\�O'vuz���4�O������)>��<>����I�>/���t>^�����by��3u���{�t���i:C{�ct�z����G�������jJ �����܍��ɸK>̓y":���	~�p>����Y��x_5��'�2���85ޗ���㸋fS�|x\-]��a6�:�Ƈ�Ҹ�<e�·��!��`��ӕ��@x`�+X0���y��j?������}F�޸��y,���
�1�<��@ei�F�=#[�=x�Z&�������x� w�ң{��C��1�{����t�U�]t�ٗG�IP#�x'_��0__5L�=Վ��'�C�r��;�=d�^��vA<X�A:�y[`h��۴I��j�<��[a\� ���:��~	܎�~�n���Ǧ��r_Cv>�V���}�yCv�V�ٽ��,�&l���s+8���҆��ܤs�5����9~�CO��О��9��yK�������g�t ���({��ѳ�-D����o�*���7�
z�]���-���pX�S!�JG���I@�\��N���.�(��w:�c.}�t�� ۊ�U����$���(��	�����q>�,#�,���y�3�2�z����-([��J^�9��Į"?{g�ӠG��+נ���.d{�V �`-��-t	N>�
�V����K��� �N����MB�^R��~�Z-�.��v�#�K#�R�A���?�K�pe6�J�2§�d��zI kM�d�V@�*�$�����4��\���G�w���!8&�����i�@�����f'o�[���L�#�d>O�+������R��b�22_]c �詮��_J��f8���
�ބ4�x"r��A�F��@71- �*��"�/�7*��N��&zD�Qǀ��Ԭ.��-��ź^�~��b]L+��~�:*�������������8�@#|�l%��t�B����4E1�GӍ�u�1�/\_���>�R�$
�t��-����7	��ն�'}�M��k$���u~K}]�X� ���Y�>��y��%K�n�ٰ�F������A_^�'?��������ō�$𚨗�*�^�[_ۄ�w����ϿoF'K�ہ]���>��+��W�⬓M~��U��|�%.�<m��էM�Ƃ��l�l�����K�x�غ#x�ط�;B_և�����{Dc=z�럱oi4�P�q^��d��ځhB�܄�������[ri���b�P��<�	/aK���d;S(Q�OI-�P,N���d'�^����� B�A��a	����_8�Z_O{�o��������M�,Wha!\��!T{
sh8�{���1�ҿJ0r��%�慓^8������ׄ�j7�l��:��֑����	<��0]����k1q�E�V"�G+�j�m�6G[���^��0:��Ôa�0m�i�y�e�u��X2��ec�c����t*�j�굍l���6�M٦nӶ����Y�Y�y=G��ϱ��s�s�s�s����Y��>�u����1~L9�ӎ����Y�Y�y%�1���Te�:U�j�j�j��N���i�~�c۴���:�
c~v�ޱ�~v�E�ᲇ~1�߀���^�fժ5��Z��?������q�]럞�@Z*۪������i�G�Ә��}���>�.�х�7�)�Q��;+��kV�.7��9\�Ќ�x�^*>��pv8��7��0V�C��h��_��=Juj�[��H[C|"J8�۞�׍��P550(��m�ij����
�a�ne��6��;u��c�������q.GA�]�Ư�@qi;1,k��(�ۧsx�f�;���U 3���l_}�a�7/y��Ig�g���!���7�Ҟ={NӨ��j�.x,a��^�W_�v�*^��7Y{�z����UMk�*�.�-t�cW��������vkӊ������`	�zA��:묃y
�y�~m`��h�K������}�F3��y�V���xoF���w8�i˖U[t��¹/�\��
��'��G�Ng��ٸ��ͻ�T����������1V��J����B�7�&�{'�e�Q)_n�6+	1+�������Q�b�"Z�9+g!��,�#��׻u�H��}��ׯ�v�a�ڡ�����;��4�ZȮ'��@�ą)��5&�U��j�YY�ٴ'����!�F�!Bɧ\�|�%/�(h%��
i@�	N��mv��T�	�_Q����O�M>��̟?s����q��~��:����fl��;����4�q&�tu�Рkh���[�cJM����a!��w�IkO[�F�pS�Έ6 �ov���lE��	�F�+���mh��:��A(�d�cc�����on�U����ӀQ��.ްa�˗�/����=�����o�j�8�Gׄ6ڹ�П��o���UЧ����F0�x��*	*$�UNFBM���ܠ�oԹE��a�%��m��]fn�^k��C��[����N���@��Մ���G���lL��S��֝B|-!�ۅ�ߎ�1P[�ԛ������@��CQpKW3�|�zZ�@��p��'�._�����ǿ=���oܦ�W���mc͝�h�����隕+7׬^�)��\�p`�;�����/�n?K��y�9�-6�!xJ�<u"�ą��HM�?ؽW��ׄi5�7�m�h�qf	�uj�RM�7���R�n������#�d���_h<�3�Z�~=Թ�3����B��}L�o����H��6�Uٰ�iP��z㿩E_������P��=V�"�vq�l٫��T�A!f�Ċ x��p�\�n}��E���[/p�| 8Tb!q���DR���ҁ�:hVd1 �\����|2E��Nnd	�5�����A�2��1�_U%*ߧ��D�tF+�����kM�Ren�>���'JG��~\?�"ݱ��zɦӔ�|��G��]cۉY���bsH��(8[4?}�l{Y�r=��Q�}�&�uU��gp]#=��RA�D�3�+�)��)/�!�%>�W�H+�O"� ��U1�h��X"�ՌB#��J"��s+b����GU-f�&_�Z�h����:��C�� j��g2�y����&N��q�V�+s]�ԋ)ܦXL��Q����'�S�Q&Ky8+����O�ӳJ�/���7(|߭t�>_��|/�|��z�hSý����X6����bm��,���`�1�h1�W[WXyF��J�1;&��'�0�aҎ1���?}����gS�v�F7�rZJ7w����8�o�o���H�[�f@�f�G�Ƶ�j,�I��F|-&k�e
�����z��ˀ%;����޹c�_+IM7�G_ ���:ɴ<:�&�G�=��]?ёt�O?�V���"�0O�c
�	� �]��w�k���Ǌ�OV�Zz�����	ޱG��$�v&�i>�!�=�P����{H�/\�|S�n��ʅ[�W"�c5|x����&���'�G�i��ʑ�Pҡ�dp\Ǡ`҆״o���vA!6үU��7DH�@�R�~�r"���ל_xߎJ��o�ү�h�0eo��{��>}������B��=���2�����������/�v���4�Ϛ�'"�UJS�A<��CL���&�Y�FTBj��4,��!�kt`�I:P���p�e�!���W�,ř�&ICx/�G�� }�/���`���K2��d<���<Yi�h�Y)��h���81s��>�Z5M��j$��04�7�bO�����;�9�k����N��jiKy[s��3��;��Y�с��y�����r��:"-B(���>�/�6�{X��Y��N�f��j��ox�[�OTC��g��V�_^�z���@k��������������h�˶l^�l�e����p�zҮ�������_� ����!�_N��E�"���~�H�o��	1[���`�
	Uh���	��ϓg����~���X�BۙH�v}z���tyF}�ؠtަP�(Z#A���D�����BM&FEd��*6��;���T���7��_��vW�3�9��X_t��77�~���������7���7��ၽ���O{�|?%q���Y������w����1��q>�at�ใT��AhM)n�R��|C�˽uIdI��J��rA�U�?�ZlY,����W.��������3Õ�"�Ҹ��<�a�5������W9�uX����@o��X5[�C�Z�m��5�3D��r���+���Ǿ�!&4��1&l;�N�����^;�lo�=p{��`��]BA��"]錄��W
�8i�A�͎y���7�/�t���p��~����r|R���U��tv�޿)�/�P�ԆŻ򦾲������ק�K���������l- ��'1q��6_�kY�z���vO��6MN� �bc�ã�p?�*��+�Ke.-�����ћo\��ѕ+]����'^���y��jkY�{�?�t��lNF6��?��'d���(9	z" � l[�}�NVo���W[�����F��`��S�}Ю���©[�JĨ�e����4�*�nIKY��;mS��=�  �=��A����{�
��� �n�E%��}V�7��O�
��?��B.B���"2<�;���P�|��W[�9_���E�]�t�UK�.���խɜ@�A��G�Oн޻���K^vӓ��=Iq���P�j�hmRm�7}%hu��ޛ;p��ni�����vm�����"��~��~`�.��vK
4f�d�ql_�񒢓������q��j�Ǘ/�kgS��^<3`���@ڊ�h�������*�_���"} 5;��jt5y�G;ae�LH�4o_� �/�#e��r%V$�8�
��z���L�>�.r�����Z�����Z��{g䮭��֦��3�x�>R�w��ȸ.A��v],�U�6��!mV�rxl��ɮ'�w	"�m����q$��K{8��2��~I��[�w� ��0��ۛ߷l���._�����SweN�>��呛JN}����ѵl����������^�o��`T���S&�A�D�t���7┐_;)�ȸ@��L��;j{{�FFy[4�� ��#t#H�/[b��B	��K3�xUmm�ݕx�l��<���i;��~&�v �%b=�F�d>Hl��O�;��T/���d����]1�q"ap>C�)��Ӓ�RZ�FCkk�i��k��6�����q�t� s[�Y�TS[MS-m93�5a�W�j*�-2�3��yҪ�U�k�i�$���b�����\@&�&�S�q߉��$6����mX�h������ɬ�U�Y*B��_T��`S��+�v5����i}���yO1M�&��EJ�Vd���s����� ����d&���O����G�����~_C2KX�����U��;#s �z�v�T��(�j�����̩c.��й���p�����ן���O���z���:�-�`�a��q]�}-��th��Z�V;��v'��&��k�����Mk8&8)�~c�~[���~Y��_"���&��)�|O7x��e��@܈%F��bL1�K�5�kX�am�<�ݰ��:Y�)��E�"�"�"�"�"��mֶ]�6hm��vkۯ�6$��/7�6A��P�,��|�v��ZV��or�=��J��3s����k#�.�4�f��������l��rqU�M<,��o ��~s��~s�~��W�F��[��8#!���F��j��&r��o"�o=4Pߦ|�㭊��_V�zݺ�k֭[s���__�y�r��K~x��[�w��aS�ҞTdYQbݣ�x%�}�w\��}��fz���=i�ܝ<vlĶƭ)��O�^�l���Kbk��W�l�ח���5g5���	����خ�N�߻�p㳈�����G�B&/N�x��Q�	�xb��_<%O ��9aZ1qvb�v?qP�_����1~q$������t�nO���x�n�*K�� �<�$qV?>7����U�}8{aX'#�^�n4�ӅT���\��+Un��9�CH�̖[�U��������~�ꈣH�;���v�O�IK�jl��e����8��ʔ�#eve�-�c�39�f�wj�ͱ�3̟��k���<8sƑ�y�~oN���˯߷K�BTԽ��G��o]��px�Ѿ}s'.��|B�/|�����%��Y}
v�+.�G5��ď�0���,�`��i����|J~����Y��ct�>eJ�۟��Gl��S������~�l�Z:ԕ��S����Vz�&�lN��q����VؘhL�:��}���/�������Mwg�����cwN�g�>��c�2�h$?�⵪������Om	�p�<��7JTURH�I�C��7�%\�u�?ta���#6fnV�E0&Ά�ix�1�D����`/��{�n�ޣr�ب_\��+��*N�^V�eM�2�
"�f��φ�m�-����5r��l�Z��o�y�H�9c;�Z�'��g]��x�uW{Y�PJ;�`�^	R�[�Y��Bm�	N����M�f
7G��~�@m���y�-ɜbI�eoζL�h+`E�@)RgZ�f�y��
���� �C�4�j��z�C�Pu�u�u�u&+R���B>WY��S�.�Bn~��Q�{���'��n�Ƀ������f	G�������-�^�C��d{\�w[o!N/f�����?���q�{�x�����N���&>�զ�~>'Z��}��������J���o���G�7~%ӄ��M�b�egf?��-Ȼ�Og�~)~)���⼫��ɇ��;?r���aQ+'o(�w�}�I�JG��������m�rJI����^e�^-$,�Y�+�2�+��~�J]�'s���GV�Ψ��.>S@>�qRJ��`i��}Z��
;E�T����۴ ���P|�tT���~I89!��E4@�m��Y���W���K��.�<\d��S���E��kkg��;����#jϞE.�������/x$䴑��$!.�n��>փf������*�-&8��˄��7��;��$KR�H��D� ��\�F�N��-��S烘5�tn��P%���9�5�ۆ�����x�Ǐ�k8iP.*��IMVgJxG}G�2�E�n�v��YB�i�s����6�7Y|,�-[,�[�Y+��y�x% �{��*l{l_z� �x_���3�g�o*��]���p��]�w�.܅�p��]�w�.܅�p��]���}����p��	��6ԧ�o�L%C�wF���5�՜�~ţ��t�5�C����׸�^�y�����'��>��9��wG���6%�pW���pW�{�+m�z�v�5��+��6�0���������ݪ���j��B�����ϭ(�QX������1}�#�����"?�$ґR��/.vd�Q�������Y�yQ����9���9�3�+9���RGy���\G^YINQ�{LfNi�cLYiYBY���+*��J�Q����c��5���Ua�ª��A��y�UUYV]��_PV1#?�4�*zv�E�E�y�s��ˣS�r�K+��lA�਑G���|�����ݢ��QVk�dМ�007J�������l-V.����������e-�X���%E�R�]�_���fT�V��E:
*�<��aH/�QU��)��(�*0�lz.*��UrA�YU��RDNnnYI9��U��^lH��5L�$���9r*+�r�r�$�[]�_Z�S%�)(*���
�r�#���j6d�MRR�_^Q�W��/�������U���f"�����<A�좪²�*SR�ZH��0D	�Օ/؉t��K��~+#=ֈkF�U8*��.�.�[,-��r!�*���B��Jn� �PP]Q���ļ2GeY���z����*�cȸ&)�-+�+|T�Z��(gz٬|ɁaE��F#(-��*�^���&0�9*s���|��@�<��e���
GIYE��vT�-�/��BQQ͟����K��
����W��� Ҝ�<ɹ!:�_9���8�B.��_Y4�T�1�xnya��$,4'H*�7=�-W2,.�XN��H\�ܴ4a���sE�L,U�o��cE�RS���"���|���ey���F_k�8�I�A;��Z�Mk5� ��UV�HX��*x�#��.�3�8_<0���)̩r�Tc~is�`�&�sT#Dt�5�+a����ʲb��RuBQ9�bA�/��9��� c��Ҳ����V���@b~q� jd�#ylZ�#slrք��$GJ�#=c���ĤDGX|&��"R�F������������Ɏ�����)i�������L��Gʘ�Ԕ$���O���6�yic��)cR��4k���B���)��I�>��	)�)Y#�)Yig2��;��3�R��K��p���H���@������U��$�	 >6}bFʈ�Y�����HGVF|bҘ��ё�±`9�!�D�J�p$��3GƧ�:R�2�2��ǈ�B:#�Ǝ2����26͑�V�R��������1����1�#�2��\�4�CL�������LO�"�cJF��,9��$R%��Ǧe&�;�^
�$� ��7\R&�O�O�،�FR&�d&E:�3R2	�cA��'f�A�Byi.z��D��ցQb���Ĥ�T �d�6֕4'7��Jض˹��(C�?#��A &<��k��&��%w#�59�ؒ#]�W�X7v##����G���Q&���J���K�\�^eN1ì�Q��9ŘV�Hfs�ro��E�2���
�đS�ފ�y���µU��@�Ғ����r�TE���Fal���$%E���J\�K��Vr��*��<�#W�rX�p$��d.� Ed)$U�A��\��X��t�p���Bb]���$���H���R���_#Tp��F\��.�|̙�:#�$���0�TcD.�� �9ҁ��� �R��3x�0΁�eX7G>k�'Sb�`T)JJy �����U&qƂ�ޤ������q�^��*���*�7H���<��Y�qe�Vȯ�s+$wQ���9�d6hy %Zr"����r�,G_��6_ғO�=�v�ƭ��u"�U�?�,��ɕa�nRC�k�%��N+r�A˓��m�*�l�����;���+<����s�VK�T@_���h��K|%[����|_3�*���$��4�q5CÆ�EJ��$��r~��+���(U�4\$���%�%i7�*IEs�ȑ_�$,�܅ݍA�6h/nf�B[aV&5�#}�!���R�q�"��̅U�H,U�[>h��k#�M+�� 诂/v.Vl���)G]�U�%�M��I���M��*�Խ�ϯ��\PV-�2�-m�PF�*�dJd�'Gn�ͬҠ�Z�0�C;�]"���u��Vbv�����g��R���w�K�͵��\�%gP[�h�U-�����R%��
no(����a�Ǌy�kDʫ��L�ȕ��1�v\슒n�ʵ�$�E.JI��r���2�t���$p{$�K��*��u�J�c��<��9ǥ��q�mk�4�H���,�;�å�y���-�̕��( pG5��/�2��H���"���&h�rE=�ǠT�4�C�V�޿�*����%G�ss�')�*�����sb�l\�Cs����^��|*�'�����r���D�/S�|��r���.��yE��+\(_�W������2�~�r�wŻ�f�-�ʓ���/�5��r���u�<������t��e�V�����YxZt����ʵ׈�� cˑ�5�q�����c
e�w�k���|iQ?o/ww���i�+���W�/�+a�t�?��J=�{v�׹=Jdō9H�kFs��Ң@=å1c_,��m���~���.�r���I��:cI��:cq�E& �̐��׮8��e��x܉?��(�/���a�'�-0�%�$.Gj�{"zn��w�1>���$��+b�L�u,���������c��/��{�AD6j��&�(�!Ǐ���f��i��T��ݔ��]��t=��_f�*qM��'�vZ#��.J㥌f�s8(J�w�w����)�\t$��M�<$��K���ЄA�p����Y�
�R�kd��P�(�UG�^���.-�v�(�,:���7��)�O8$�Y�ɒ��~7^�판�4��8�_���X�B�|&�(��82�C+å����r�x)��;r���\;w��
#$IRR�rt&�$�<��c�c��u�K�N���H���pɣ��X5�eS�Rv͹0<D��ą��xW=�CfM�Osiwx���J+�]*�/&�Q�Rי�RH��;�E�8s�q��>�6R�\�n?r��wb��˽vs&J{JuQ��(�_�kĮ$�k��c�k"�5߹=�Ǧ��3��$M��30��9��Ÿ�^#>{Vә�3�����>%9}S���>��m��<��<���`ecVb�e���l��iO7N�%r��y�R�kpV����_��lA�Vyi����X.�{c�ٲ]��Lծ��^�SqE�Sկ���˯ɿB껜g�")a�OF��V���I&Bƻ��Zo�>�mi��
��<ϥq㽚X�j�>��q>$���N�OĈ���@2�EI|��nW�l�l9ی���'��h�`�G{'ۍ��l�`ϡ���G�O�%���h��^E�5��g���*�	UT��,W�F��r��;h��|��g^�*���y]�=G�m��E�l��1�R!�w	z�d?��h�ɩY�sNE�t�;����Q�� I/�)s���9U�8�*RN��F�I	Y	��H�Cu�в���Y�!��1�g��Se=fl*�4���I��љ��=��T�Q(q�:R�}J(y�����'�qH��*9ԈIri����lCBHg�MzCaZ��B��/kd��s�C\��t�qoyи�>eH���v��}o��/D�H<�k{�D��٤(+o�"f+��z����X���3sc0ZЎ9,�&j�S��O���R\��PY�,��)�M���`��_��XO5�%�P� &3�'���HXq���A�
�SpO��x��qb5����/��\�1��G{v��(u44��rNC����0�s'z�p6�Q"9|HY��PJɳ67��~���e�)����o�Tg
�2;k�ڳ0֕E�>l�c�,�e�l6�屙���b��៏����l���Zv��b����=���}Ů��'\�6��y�Ļ�ޏ�	|$O�Y�>>��b^�����#|%_�7�|�����!~�����w��c~�ͯ�^a�Y�Q�`štV"�Xe�2TITF)��xe�2])TJ�*e����Z���IyJ٩�Q�+�#�	��rQ��|�|��)�*?*���Vծ�Q۫ajW5J�R��d5U�P��)j�:S-Wg��������u��KݫPkգ�)�u����������zM���҈�i6�_�B�NZw-F����Z���ݧM�
�b�B��=�=����i���m��O{A;��^��i�hhkW�����M���Lf��)�lr�:�"M�����D�(S�i�i2t�-5���	��"{P�����
c���*g�����m5�G=��E�f烲^-�7|*�:�!�v�XaW�#�Q�f9�Q;���:�m��6M�v&��'���yh�6Ґ��8�
��S�� j����O�W�G�����w�T�͖�H9&JD���������Sx{���9����A9+j؍:Y�.7�KeO���dϽ�Ζ=�d� {���a�9U֓�O��ϹU�EO��'Ȟ,Y#��z��_Ԡr��q�oȧ�EM?u@�\�F�tYWIJ&����E�Ȗu��)�q�ș-k�@�3试R2���<9�TS?�q��T�*�Ȧ�A������5��m��S��&����!1Yǎ �� �9Y:I{�ڗֵ�h녨��:Q_-)u��$+F�u��Va��Hi<��?Rb){��U�Iú��,}Ǧ7��a����h�Ӱ�;��H���/7��6�r���RnX�J)��:�A-z`c�Q���Z�_��T���1^5�.�<��������Grּ���O��A����un��F�Sj��O9�ў�\,��A�nx	� ���g����s�y��J��;��K��_�s$�er<�q�s�.r�dgk��.r�8�'N���S���X����O�������x�p��pu������?
^�� }���#�`sd43bN��CzC���q&IDZX�VWQ�oe�2I�$���(ϐ0d����-�A�l]m=H���=d�-�6�̱%���y���@?���B����ݍ\���I��OvzW.��/�2[5�����-z&��Z�<i�ٔ�h�2z�n������g���&{�r2�2c{XY�<�,E�.~X|ۨ�>M�=���ͤ�CG��?t;�4��n����S���`zЄ,��[��9}��������
��^�7i=c��|X f֙E�X6�e�lKg��d6��RV��E�Q����mbOᬲ����;�s�[�"��>e_�:�-���\�Vn�mx{ƻ�(އ�q<����ͧ�<>���Y�A�0_�������{�^ˏ�S�u~���?���5~��R��)6�_	TB�NJw%F�V��J���ܧLS
�b�B�+zDY��S6*[��ne��rH9����S�Q>P>V�(_+ו�J��T�����C�F��� u����R����du�Z���U�<u����Z���I}Jݩ�Q���#�	����zQ��~�~�֩ߪ?���hVͮ���kaZW-J���d-U�в�)Z�6S+�fijk˵Ǵ�m��K۫�j���)�u���������vM���2�f��&E��<����U���R+���ݍՋ�lG� ����h�����"�#E���؅��"sP�,�I66�_G�#�if�G�x�V+�6�vQDr����":)Y��UA�V�G�_W�#�u�)I���""�u��Uq�*��S�@��T���}�fS�t�q�%�z�G�T�q���'�z��d=M�~Y��'��Pߧ���;�)�s��ɒu�򹈁���S�����T�� 冐�'v�0+W����w������JJ�e���w�����7�,£�UY�����~V���2t�Q�I��7�*�B���]ɩ���oY�&������]�,e�����m��s�3��!����~iu6��[��b�X�����(�H�H{.,$R{\�Z �K��5����3Ѷ�3���J+�m�=C�"4���m�V�r]b{�C͓�4ii����i���i���G��v�3"&�e���i�"�@�C`�����l�^I���,$�~؛�F^�"�� �P�K;��[\�/�������Vi�T���H����E>�W�DH���D�Á�v8�yE�\:	�"�*������G�?��+�o��}]H����#��z��@O��r?�>��H~EF�H������a?*�����b���'���4墤�^�`�,�M�M���ǪH�
�����<�����B�s��d��q�W���2�!4� #B������4X,���s2\�"[^��û��^̢���`*�~K˙8�t�)��i��2�˿6�A���"�L���+���܇f22�<�<M�q�~�t��LW����|�P�3Ŷ��xRbKD&�d2a��]��|,�Od>���������t'6��Y�ĺ�֏f	l$KcY�>6��bV�氇�#l%[�6��l�����{F�*;��a����5��n�z.� �����;�H��<����|<�̧�B^ʫ�<��?�W���M�)������A~���g�[�"��?�_�:�-��늢X��Fi��)]�(��2H�S��T%C�V�(y�L�\�9>�,WS6([���.e�r@�U�*��ו��{�G���W�5�rK%���T5PQ;�����:XMPG�ij�z�:M-P��
u������R]�nT��;���>���z\}U=���~�~�^Q�V��7�z�if�GЂ5��Y��b��P-Q��k���t�P+ժ�y�"�Qm��[m����Sۣ��jG���-�vY�T�R�Ӿ�~�t�b���6���0SWS���i�)ΔlJ5e��MSLy���r�,dq���3m0m1m7�2�50՚��N�^7�7�g�����+�5��-31kf���h1w2w7ǘ����#�ifD%�#�~^�t�lϓ�-��'�{��=��F��s�i���n��m5_�c�W=z�{�gyb����Ǻ/��ظ�Ei'۞c�������V�D�1˓�_�ޡ�9�~-e����}<p���K��׿���T��tJ�z֞2t���G}���Z��՞��ѿ���d]?�6l��&9x��ciH̞���9�n۰%me`K��z\6�j���ϑ�7��Y�imD	�=-�Sz����k���U���K�{�Q4L��m6�F���Y��=���)������Z�4�D������Y<��i!���#�H��3��ӡ�;��Y�'��a���!+�&2�l!ϐ��Ԓ	�9A
�)r���3�ߐ��_H��|�9#�Ĝo�w�	r��@j�-RO6'��Vj���Nچ�%��`J�D������WuT���^���{��GB��4R�)B�a(���)�)bc!PBӀ!�1R���)F1��ƔB�4����V[Ld#bDDDDϞ���>^&)��d~{9w���{���{wOr��?�~̳�S��o�������K�R'���\R��[xHmS�xXݡ��)j��.���︈����7Wږ��J�:�Ii�8k�io� �y�\!Wɵ�2y�\'����&�En���v�C�+�ɝ�1���%w����5%�DS��e�2R��W&)�J����+EJ��@Y�T+K���*Ɣ5�uJ��Q٤lU�+��7�}��m�r\9��Q�)�+���I�dD2##"�"Y�	�ɑi����E
ňy�rD%�&�4�"��E�"͈͈m���ݑ=���AZ[�(�m4r6r>r	�W�J�ᨎp����ѡQ��Fq��ng�Q��(�p���Y��h��;�6�@T!�/�.C�D�!��M�D+�ю�����!D'��$�+����ˈk��aDT51�E}*z�:11�#�:1	���Q��|�H-E� �����v�.G�RQ+�:*=H݈؄؊؎؅�Xݧ�<ؓ�G��S���z�� ��:�i�!�C&��Qx�^&�dL�!f �P�P�E�?S�G����V�Zh���;@��N؍�ʇ����pN�Y���;@�i�;u�隫�k�5|;�����Ps�x7a�m��o&�zZ!����PsZ�G�i�4ԜVG����Z�֢�j�3u�u �"Po�MC�i�7��u!�5Ԝv��G��;{e����tԝ���Qw:�NG����Iz������z�^�/����}��J_������&}��]ߥ�����o�G���)��~N��_1��� �6Ҍ#�a�2��	�dc�1Øi��<�ܨ4j���
c���h06��fc����m�1�2����	�q�8o\2���������`s�y�9�gN4����\s�Yh����
�ʬ5��+�:��\o6�-f��f���^s�y��4��'�.�ۼ`^6�Ya+j��o��Xì��k�5�ʶr�<+�*�J��"��Zb-�VYk�uV����dm��[��7�}��m�u�:e���Y�+6���`�v��ag�#�Qv�=��lO�g�3��؞g�ەv���^a��������lo�wڻ�=�[�A��}�>a������K�UGrGw\'��u�uF;㜉�g����r
�g�S�T9��2g�S��;�&��iuڜv�����w9��1���t;���57�F]��݁�w�;��w'��ncn"Q�@�u�{]�^��E�u�{]�U]�_��E�u�{]�^��E�u�{]�^w��E�u�{����g���.z����{�Ş�y^�7��ey���4o�7�+���y^�W��xK��jo���m���6o�������{G��i�w޻�]�%_�u��Ӆ?��C�{���8�?ş�����B�ğ�W�U~���_�����z��o�[�6��������C~��?�w�����-5�M5S�ԁ�CR��F��wߛ��YQ��|��xl��D�)6� ��c��������`;卵^����������s#��y5ɫ��rb�<8'#y����G'��g+?��x/}(?Y]����]��>�Q�ߛ4��^���Z�aG�����纒�AK��-1�|�ܛ4+�Fvի�s�6�5}}W���m�+��D_뽵��-�b�C�[)Oc O�gcm��<�Ǔɓi*(�}�lbpw����٬��a�6��ڹ���A���#��UA�ldI�' ��<��"0"G���S��60���J��+$	���یډ�XoF�d�[��$��{y������֐�'�g�����	���|���L�{�}ے�X�8����#>���l�	��D���F�S�����２�T&�y��t����	:z�����xE���R9I�$�By�$<�q�g��ت$�۴'QG�N����]���=Ϛz�M%^�EV��L6C#>�����q����.��'��S� o!yK�<����?�,����C&��I׶o%��L|p��O$�N�ӓ�9��zl�m�bW�x �N��5ݑ(ORW��؞Jݝr^�tGϊ�~ҳ�L�Ø/�=y��?L�a�Eċ�W�$���Zi���	��� � ���g/#^�c9A>��T�����Y��0��e6IJS���R�cI>�����7���%^L�8��_���<�we��z���8���X��e�ˈ�Gy�rQ��h�g4ֳ-?�b�4�d�e�����lkd��'������g��v��з��K�)�2Ry������?�(i|�dH+y�>^�(M�%�i�����O��ZëC���u��C�|MJjJ*_��?�����R��-)�Rv�W��T�I���������|�\/��[���o�Ղ�[�V�M}]m�m�Z��Vv��UO�vm�6�w�}���(^˦H���k�6�A�YC(.��Ⱥ�vu���b��8B��A�C\D\a�0!�}6"���>E���Q��	��8��C3bGO��ׄ�1���8,V�9_*v� V#����q�,�!���K�݈=���AZI�\��:�u�F�E�gw�;�Ҙ���o-SX���ok+?F[V�Q����=R�M&�S6�k�2��ձz��&��ZYkg�G��!�Ɏ����u�]f�x�G��}>����H>���x6��y<��R��/��|	_�W�5|o��&����;���}�ɹ�u�y_������w���Kx����E\2���{H&����7��oV����z*�(���"�!D���X�����~X�3�Oc-���*��)]H�o�7�����x���G�q��)�3��>K(�>kќ�E~���,�����7#5c���m$(c�L}����Y�Ï�b:��L).���B(.���B�Q\hŅΣ���-��Bt?����x$�$b?㭐Xt���s��9s�^Ħ���=ɦ�+���r�*ʪ�,�f���㝋t��sK�XE��YE5лx����}��J��`7��8ł���,��?6��c�شx���xI��C㿋=�b��L�(zz:vcyx����ձ�_�뤸^%S��R.�H]6��Lʝo��rأ7�@D/��؇��$���c�ɯI?��g�>L�uI�/�_R���|��ȩ<QN$^v��C�sC�mS>/�	�h�El,����<��'�1�$|
����l�OB<O����Ex�������-x�/���
l����Կ�P���C�D 4� <�?�>w�p���=��W⌶?E�ܥ��F��Eb3��0������́����/���+�5�<߆����=�>�
w���տ�T���S�+� ��z� ��#�k�0�}@�(\�Y.E?,��"b��Zl���������4�vdC��,(�"(�
��j����V�jX�� ��Ͱ	��6��zA�RϪ��s�~���^�t�k���e�A�A;�v&�#�~g��"�z"W&ك�\؉g��> m������:��y��t�(�����1�٨��G����wݴ\	�ϐ6R�Ų�������w���_��o�7c���^���
endstream
endobj
30 0 obj
<<
/Filter /FlateDecode
/Length 463
>>
stream
H�\�_k�@ſ�}�>��7� ��B�[6���$+4*�o�q��+$r��w\�z�����w?u��i{���w���<�Ă��[���ݥ��������~<M��Q�;<�.�NO�tt?���{��L�CЇ�<��*���w�p�[;�l/��h{��������{��}v$��1��:����xv�+�UѮ	WEn��{�7�Oݿ��qY�7Q�[���3����B�Ba�l�0�8L�@1����KXA��`�0����-@	P��OP00p%\	W����00pe��%a��� �*���Z��kU0@(�ת�yu���QMZ�<�NH��Ma8�0"�02�0�P�#��&�Duf��e���`D�]�v5 ���cZ4�l�	$�$�H$��C�����eJ[��պ�_;�ݼ�?qO�F����yu�ߧ  ��%
endstream
endobj
35 0 obj
<<
/Filter /FlateDecode
/Length 15605
/Length1 32980
/Type /Stream
>>
stream
x��xT��?��^{�=���FH ��$��D�	$@ $!	��d2!�$r!D@@�*F�R�T�Rj�Uj������Z�V���O�kk�J�m�"�=��ޓLh�w��眇,��k�˻�����0C(!ĉ�L\3fT�m}��g�l�Ao�̂�c�N;AȆ)x.�YVZ�}ލ�̈́H��Y1���e!���+J+rƝ{�ӿ���/�6z�O++W;���]��z��'i��0���敍�<��S�݇�w���6#
�0϶���g���-!I�'d��:���|+ً�Y���iR�k�<���m��{�b\�c����c�ڻ�����Y�^����;1���i�=$�=@�-�����om�%�`;on�5O
l�DH<���^I�z~d.6-���9I4������_��E�W@�$��?XglT��[�_V�*I�$�?2�c�E�&�%b'n�	փ}�-z/QQr���p~�wH�����̘l��O�!PN:���.������]��!J���������}���[�N��J[iy�I$I�s����]� �"��Z���z�?O���� S)F1��|�EbIk�"����'>��$�"���\TV�#e�eR�BN.Q䷓���/�z#�C:H55�UIn�N����?�n���,i%'�Fr�,	�%%�Grb���V���Nr��z��Of3�#=4�\�(MŪ��er�.�x9��;�+�����L�Jࢠ!Xv�pP����l"p�+��@E�^n�K���TaύZ	�����N��}OhU���+j	8R1�58��W��|q����"YL6�:1�>"U�����OF�r`�)�A6P��q�.��/x�K�_6^��C7NB�=4C�����w���ǐ��rle-����3[�L�Nf��db�=�>�6Ix�-���Qh�#fha�Q�j#�E���d_���d.������t~�g	�,��9�|H[�cd-m����^�f]N~HY��� ,�wH���'9}RJ,(� W5����!��d����x��!T���th>	�M#�֡<�<p�>����;p  ���4����d�N�_���~Ka��d�$�����$t�h,o�]Dބ\��$��ϲ������|��$]�w�;�������s�������C��x4�9Cn#�O
M'*�O������n[A�:��E��k~@�!��;�e�F\t�&��9z+��.���e�}�~�~&�J�t�Aߡ�a��I��Nߣ��w�B?���g�z�|B�=���C����~�G�G�=�}Q�
(���W��ы�������3t/�1�9U찙���Iw�l�@@��Z:��QYN^��<B�A���ɧ�$�r�K��)�5��������O�7�1ER/����A�N�j�k�O����.�r�����$N=>w	�[x�L\���	?� ��x�ړ{��&��sл��ݷ�څka�w��r�v�d;�6�I�����v��S��_0ކ(�'V������$��o��z�<In'���g��ж�$6�s�/c�#�����S���->�Ы�"Z,��&�9�>�Ă�(A��w[�<�]C�NXJ��/X���_�{��/��π��� @������M���.���gz�GI&�oM��*��Q��VPzW������a'���,t��4�6�
1w����4`�	u�؅߇t�������R	��l}&_M����=����;�}p�c�n�*��ϫkJV�����_���-̭�7/�7�SL܁/����Sb
�	��FTr���g���'AS�B��QR�h0ϓ_�,�.'fX�c���A)^k/��H��}�B��Ix�2<�c��>X8�CZ��[Y�G!�����ȿ������7. �r�V��%�E�;��i�&�Zϓ!X��=�}:Z��w�F^~<֞�?�����t
ZB��!���x$�.�do!�О�'Y��4`�2� '���R����EX���o�堲��L[I<����o���S��S&�	���(_���p�)����ȯ�_�_)2br���tM�4�]:�2�JG�N:�Z�M2�iƋ��h�i�/���[0�l>����t4V��~3֎����C�g�ȿ��Bo!_b�p�JT�������&�2j&h��9���`�EP� Y~σ4yl�Y�����<D�S��Σ�������*�b	4���?�jh&r	{p]���`��j�Us�:�<�2ȊG'����Q�-��ˣ���� �=ʖ��i�z0�s�#���ͳ�Ъ�AZ-Xx�>�~X��۰�8����J�9j=����7p���ާ{?Q�@| �v�L��Px�K��D��k��e!9)2�j t?��2�<���P��k.���.��x�A�h��[b�7�x��2���h�е"��;Q�Ù@���oD$5#�^�yG�VD,j܁�;�}<HE����������8���S�HXɱBvPC���	���S!2�7�kR<�����f ���穁c�|i��.�ސ&�G�z�\s۞�.�D.��LENL�k�����GMe���%��s��x�ldB#�]Y��	�%����L�w���O3��YX���"�v�N����JD��c��ϝ���0+�1��EH�
ߘ�e�a���e�"��1^�v�I/k�/�r���2����Q)F���L�G���Z�B���^�FB�xO<�4�MC�4��U��5q'���w �![Pnׯ�ȃ(�_;r�L:~����B8-�l�_/[@��y���*Dх�Y��e��l~:P
<-U+Cz��AOW�;P��e(��JY_�2A����B߫�A<j,�����!����Q�A��cR*	��wĀ҃\d&��x�(<C�7Bg��U��y���ls�{SCF<i�u?1Ή~����	b�*ޡ��:z9Ff��G�� C���W9�x1�!��I_�8�=D��F�W�dE��8b��9i}'�)�wi��W��6�������U�x��u�����^�}e������1��}��N�����^�s��:"�4\���¥[ o9���~�>^گ
�@'҉��y���S��~��'�J��M��s�>�h��ȗ�q��L��3�����'�U��~����oqzO ��H݆��1����B��GB�/�iU��v�{%Kǒ��g(w�+q�-^$G�k���\dr�q�_��%��S�<�!B��ѯR�z���'_�\�V��sMZ�5���G�2�>���3��x�<�s�>�.z�(ɡJv�iI��a(��6�.]��t+��.,SP��Z�ڂ��x7L�A3���]�ɽ�]2�,���#��ϋ��*q��g���'Om?e����r)��dk1����]"�5,���&���~a�p� �[b�NO�^9}#Q3P���ԗ��ߋ�w��Q��|��#PQ��uŨ��9�娕�P=���
PP��y-�m��Qעv�.B����C�v��<�	*�q���|�V2����U���!h������s����i�S��X�)4��=���-�	��K��S �̀��f�Y,zy<��U�{9?����X�Z:�y��"3�,����ZTs�=���ʢ��Y�]v��);���	ʪ�xe�!%�K5�SS>�������U��WX�C-\Q���*4���_X0��H������?�쬓�^e��w����><S9�����~;�����Feo��p���~���T�+�����6�UvJe'Ǳϰ6���߭W������)��͞�,{.M9��s�ϥ�g��Q��Ğ�aGU��q�'��b;�����Ӹ��r��3�ϟ�Q~��=U�~��CO�+�T�d<{Be?]�W�O�a���~���~�dT�����U�?�=��=�h���`�U�A4۷���c���<�}��yȢ�Q�C�[e�Sكʃ	�1l�ʾ��=�������S�Sٽ*�S�Uv��v��n�݅��T��0��*_�~��ic]S���m�3�6�m��Re�3l�f�[w�*�Zʾ��He��l�.��6��6�nS�F�m�a�kح����֩�CekU֮���p�mkg-N��١�ɚ̯�&�5��au��P�V��+���*;���:��µa��-�j���j���yw�jp�:�yV<�xT�b�Re�3l�fy�-���l�[^���*[��%ϰ[R�b�X�YYh��g����l���WY��*�J���l���TV���4����UY�:6g�Fe��fodE�l�.6Se*���i�X�{��?����V���ԛ��2u4���nR��ݨ���J�.6y�Her�4�MT�*�p����l��ƪl��r2�JN8ˮa�_aYxȊb�V6JeQl�����J�.�����8%u���%�,	#Ic�+�%Wk��p6,���,,�-��R���(��)q�ؐ�Te��bM1Jl*�QY�ʢ�,��*s�|�� ���X6�PY8�+�q,Le6�Y1׺�YTf��L1�(�G�V�*S�T�c2ȣ�3)�QbQ��cF{h��4��������^"������P�3x����ۑ%��s�e��M^ƵJNBf�O��u9�,yL�]O6I��:�qҩ%���1��I�N��q�{�F~� ��a�p_$��$v�!����8(�D�K��e7�M�@��*��`��R&`���T+g�9���Q>C���Ô3�(c
}[Ps�>Ks��VI��%l��"w�OI���V �}S9C��)��PK;���л=�(�C^A�ȧ�"��ɋ�FBK�J�Rk1{��v���%�.���$�Βg���[/��G�2�M /�*�������he�����Md��.�J_?+@fQ�Γ��0p!ƍ�� i���]r��9��u�d�;�L+��LrN�>7��O�;}nL�#ɑ��H����V�O�.c���2�D��AN
���
�/�y&b�ل��`.L97nu���6=��ʙ�3R&���v�����ę{�;�PGV�-�0¬�p��˧&OvN����PuD9cSҤ	v);����)�JgS������}�����}�9�w͑�h�p���\�� u��J��:��9�:�K�1�h;a��9�zY�'͒�4�~��ȳ���o��X�+O>(͡����?��%B���9�ӿC��I�L�$�~!ݱ�q��vC��qGKvFE���H��$�H|����X�snr�]����i.K�_�r���F�|$���V2��	w3�:ӽ��o������ё�c H��0���9���/�qߟ�SL���r�%ǐc�1�s,9�RRJK�RV*�*��Rc���\j)�v�n�-u�n�[�6t�M��nK�u/�K�J{�^y��װ׸״׼ײ�:�Z'��q�8;.W�������[�[�,�K��r��DGR��h�d�h8�;'�L�O��0���i)��A�����M�XZ2ib�tOke���|�e���v�<�{W���¥ի˾=fƒ����ee'�������o��
4~�cǶ/�ڱr�����v�U��.u�s;���
�%�m赅T�G�M�Q�5(R�ʒW�g$^��`����	C����S���Ɏ���d!�q���2vܢ�I����\�{����})t�k�J'$]~���^�3�ҙ�!r-dO��#ht��E�3Sd4K�f��'c+l�v�J�B�#�X�N�L�����)L.c��(�A�7T��W�h�����A��p"0R����rS��.�mnYr����<��xfy��<H�)��ז��^���N<��+G=�p��~� ��d�;�Dz�-�k¼�ą�5	����i�3bq�5�#Y\d�9���b9�����\o�8o??yN��HRrZ���@�`�I'j��K�Z6�?S������[�U�����s�~���-�'֤�?Q����������ǩ������w�;��P�|�ȣI���ޛ�q��T��꾙�0�W�¬��l�(f��(�Ȋ,)�"��o�
e��V�d�ɨ�6�Y������q�NW�ǧ�!�>�0�-�"���d3M��e����4����g�|z��/�x��w�E�5��/��W�К�O���s���Bֺ�	��"q�h��Ya*U,����@�襝�\1��q�2[�է4��@A�ul�z+m��X���� }�/���{��2��%�ĥL�U]�s3<�b���v��tQ��tY�͢8]j7�8ⵘ��y�k�5��,�J�X�q��Sq&���8�+	�SמX��s�	��c3�w���Y��>V]�RR�4���Ai��='��^_u�?�oT��3���g�ƭ��{������ؿ�V�Uo�oӲ�{w�~3*����^�6�
;xv�Hƹ�7��	^f��>�k�0�+�N"��".�`��5G����T��	p�7��b��i���١ʟ���޻[VS�e��p�S����u����tՄ�j������7���ԛ�U�W7����M"~�w.��࿕T�ǘ+�B]�2*S����CD�ʷZLV��(��&��Vx�#��}�ܧ`/|�+�b�I����ޖ:�X����Au��ޏ
|��>fR��2)fb>f�c�����ȷ�L:.���2 �oD%�nb���%�W�Cw�Ƒ�u�w����z�� wn��A2RFHɩ�?#/5�$�4��d/���\㍀G�LOK�Ibd�31�0��M���c�%��>�����xo��(ax�p�92eb{u���2ɕ�l�j��흛��=��񂬒��)�WАZ|v8ݽ��4��ů�۟��K�b��=��W���hj
�~ ��"�|V�}�{�	a�����A��5�-�P���W���� b��A�=��̊�	�?�w85G1��+%��'�M�4po����Z)c�k�{�����v��w�Ts)Sz�w����A.��dY1[��9�"4T���&��B���Tl0��K�z�0�D���ԗާyI�O$���/A��t�E۷�Z��B&�����?���()2��t��@-������Md�k~���[I�}�-�^ `��aw�5KH%�dd���歭���b˳%FL�l�*F�f�a�f.	�ʄ���$!Dqn7�P|Bꫢj�E�O�K�iQF�T��b���h�DR;��v�n�4ڍ1��f�R�42)�&�3Ma4�O4��>L����RI-�� G!E�t�R��s�O,����%��a�[�S�eF��)"�RpX�-�`�6�)ވ`�n��
��u��M��T.��LN�U�VC4j�0(KA�0�B�����~R}/@ԋ��P�|�+�~)S~��\[I9|�&��C��A��fo�'�7�猈.l�\0��ze�*����VOn��o��%�M���)^R/�{t���U����z�W'�j��G����jݱ�;Y{��޹��7u"������\��>�Y$I �s�s����eX�,3�����bhl4�	4>J	��d��h�9�6�*ˎ�Bł\7�fc�p���a"�����?�|��|�9�����~q��1��"SȦ�\ Z��Ȓ:k�����jl:��5�hߛ��fԾ�����^_�3��v��ݮ������LZ�{�'�4������CV����0�nuOn2KF�#1qx��:<Q�����:��F��z���-��x#%��p�3y����ܜ��>�
�h�zj��UlJ:I��RFdFTFtF�D��Z�X��,R��q�H2���R#S�R�Sc&�ItA䂨�b"aZT�Йī�94�NO�.y}��'���7�[:��zX���՚��W��F�V_�N:�ZʞVy��)�7ͬ�>�G[���m��
��*_������=7R�u���&@g���.+" 0���#FYAĥF�}��/��?�\�d#�ǃD_�ے�� �5�B&\�3J���Y��Ty=2�l�ۓ�J>LINP"���x~�47�U2۔���H��@�]��ϳ�IBj�P��lj�J[�zgrWƶ(�P�f�&���l������,�16�ޗ:�g���2���<Xs"!!KW�~��B��ҹ�o�0bL꘴	���>�O�����l��~8d_ܾ���#��t����=w`��'ӭ\�"�k�}��R&
�0a���\x�+3�;�2�WV=�N���=�Y����:����I�m�^��4�Xt�M���__T�=�ˌ��-��~��S���Kn��������4�p#�_i�}s���a�H�2"�b����p��Q]��$%eDJT��DG�2bDJ^�����I�p_��w%'��"�R�#�!#����A�]�R2������厳��MLg��V ݘBs���;��N��*���[�ܼ�v���Y��n�ޚ<��4痛/X���͛�T-�Կ~++�\�����Z7-���߇A���k���d�;!b�}q$Y��8��Evٶt�	�]�p������M����߂��E?Z���W߲������N�{~��)��n�s��*r�3>��whb��:3�H����]w�}7O�|:�ןB��H�1sqC�����(�8G�1"UJq*Q�Qy�N3�J1w��l��+:2*&����5D�2X��qS��k���W��.�@������by7q +�'��e����7�������o������ѧ�
缶�s?{���jݼyq��OZ�m��ynG��>�M�֮[����窕7"_H#K��d{�eaڢ�����]1��|��p<p%�Y�1�e��C����c!��c�C��u�$?�S��g~�?�?��O����O}*G�ςI�=h�oo[�Z��^������nUū�G߷�.�5v�z�E��b_�����23����ո`�O����G�u��I�ݡ	��=�7��rO6(v����V��H�#"�y���L����n�a	��Y��v~8W�)��(b��R�H8b�z"��|e�'2Q#�	0���	��K���Q�t�Pu��=��3�h�=�gQ߫�y�/簷�K^�!��,���}�}0afEɎȦC��Dd'�\�p/���Gd��CƨL62���K�p�2��1q����4�k����ޑ3ڐ0,+BζY�Sr�������)�Q���s�d���t���_�Kx�HrJ_$�:Hбs%R�5{����o�H����]�wNj��˾�?uH�M���͚��������W.�`U�V��@GW���$����w�}�-���E#W5o���.�1���,�z(��]n����M	R^
��G�va��5�'�Ј��0'Ol��f�+���#�G�_��N��iD��oc�TL�����n�`P$���#�z[�����E���7=��������y����V�H�l��ef���G��2D���T�w�k��-7�΁^3�{�{"��fSl6���H5���{-��d�A�n�e��Cx���lisY�9Y�Oq���t�㧹�������rj�;�h��M�h���E�{F��+.�tw�i��O�����2$���s�?%���� R��D�۝݆�&�3�D�"�D�f��n�g?~��SszRq��9�@��X,�Ǎ����i���Te4.����7�c��m��0z�>�r��h֞Mw$�e����Bwv��2�i�oXB��8e�%:&:V���FXS�6~����%595EINN�Km�-$m��2�ٕ���ؑc�<$65�l�Y1���a!)�DKjT2I��dq�;���|��)�;�x��)�/�L��SΏ���O�!��4�9d��z�d�C�Pܓ'-�}.j���s�ZD9��q��M�mtFf�Ω�����HG����Fo|��c�Y~��%�|AQ��\��!mY�>d�-��n��x��ޔ��i�&yŊ)S�����]F����厫�e������� n]�.�\��.��q]�,���V)��3#/���E8�x�f��n�F0��Ϯ4Yr�x�t�OKɼ4_)����u����g�������|N���}��zq�����l��7����q��w_��k��i�Uu�\<"��t�KRG���d�+�'�ذ$����pF2;Q$&�A�I2�SȰ�.ǰ.�6����v�Ѵ~,j�2d6`x6OҜZ��Ƽ�>0����80לxE2JS�=ttO�M��<�T�9���f�_�m=v��Z��4��}�`�.���3��Mko���h��O�lڴ�����[yL8�;	>8��4��&0q�R̦p�#�����<T�8�7|�y�Vk�F��erB�~��B'�S����������+��Q����V���9�L��֑�3+�O/��+�xw�m�)$�{p� �w�&Eؔ$�Ɍ�˪��\yV�+I�!�b�}1ºܕ����&�p�N0F�#F]�0mW?�y�s�i:x�K�WDE!�����$�4=:=f2�L�H-�.�YD�EҢ�zRO���N�I;��趘��� ��������Ę��t�¹�Es�sb&�	t&�I��F��/x���O�!y��������'�������}/�8��M����C��e?����)�e��Nj���y���9�K�'ɒ3q����OI96aB��x�9�6�<�j�z:P�<L�H��M�!qC�7�*\����d^��}^�b�f�I,�a�34nHt�Uf�S��1Ԏx����.L9unܕ�(��<	�J\�d�&��uY��PR����}��C=�@3oVVOt���3m�N�ڸ�iE7�Y���rL^Ad�;�%�yI�m���_�h!�<�����\&F��_k�;n�/�I�̍�8Yyj7������س_��~W��`?��{�5����7�����o���&�dL&#��Fl�Ög�g11�a5���S���Q�C�@����{��u@m�%��D�(�lK��m��~e�e�����I��Xdk�)�:�����֙�tS�u1[l���f��:�����)��v�������*;M��GM�Y�Y���W��FS����G��UϫC8E}� ��!M�=ƶ�O���'�����
~E���38�D`K˜I�$ґdw~s:�#��I�5�#"y���x�3bG�Sdb4G��"MH�����13�=��٧}�\�F�Z���N��7�|膼�x`Xü�)�g�8��uZ��i�oEųw/]S)�\~�-��]TC�>A~�`9?s���$s�}��E�v�&��a?��vD�V�9Fr�o�(]ҽ2�+ʲ�n��G1G\L���tF�m �&[��ue��%����X=��8u���W?q̵C`LI�bL��#2eb�8�� I�=����~��.�b��z��:�e�8���@��>�Vߙ���"�lwϑy~�x~mV"��z٤DF"Ew���3<�)GX��e+�a�=&���#�(����D��1��xj ��>[������_�IS#O�H����C��ۜ@�1L=�G�!��s���M����RR��<��Q����C+����]��i�,�̖�U�Jy@��)�݆�x16�,&������e����r�:�zĖm�]��a��]�~<�xDL�	�H������e���r�\/���r�\/���r�\/���r�\/���r�\/!�cg���">!���}��r�J�x��1��O���/��b#z�@b�z��/���m�[�z;̼����'�����x:fY��)qYs��D­��6#c��吶B�X��mɲv�mI�>���$�����L��������tsgK�ʺ6�Ho�kܘ1���N״��ֶ��1�U���v�74����VW���ײ�W�m)��,hwy�<M+}�.O��U��jn�n���j�������
OS�k����*��v�_Kk���5.;w�6�O�3F�3����&l�T��ښ�rrjп�=��������[V���|m9���s�j|벛�s�뽾�V���cƩ��5���sU��ٮ���l��1p��4�}ܳ������gנ�끢���S�k���v�kC�X�|-������]�k�a��-��6_M����c��\m~������`����7��.^ �g���tAx�^c3��	mu�ޠq�52Y�$9�j\��V��ރ��Ao{�������o �Gr�b���_���'gLZ|�-��v�O���a���m>�ÀY������c�Q�V�oo2���F|~��J�mo�|NN���'��m��
�#���oq�� ̮�:�����l3gt��:�QG����\��-M��'��]��,Wk{�*����h<n�Jr�����zNGk��R�!O��OP�i�@�O	��mC��˥�ܯژ�����}:׀��3�N�����o�]�lW[g��փ��5��6z:9�FM}m=W4OCT ����5�q�� ��O�ب��Z��I��������/���H+_ħu�N���h�4� D_ĥ"Plj�t�Pu�����n ��F+g&�M�D|�;�F@����Օ�g��|���+��n�`��{'�k�P�!N�Z}b�um����&�n���~@$�:O����
����|�v�^�j����J�W�5
�N���n�Bt\PW� ����f�w�g%�-�����X������Z�ԬB׌ҒJWE�ʅ�兮�
WYy邢��Wr~���\�*g�ίtaFy~I�"W�W~�"ל���,WaUYyaE����U4����}E%Ӌ���tMú��JWq�ܢJ �,KuPE�������?����rQ�kFQe	�9@�]e��E��痻�旗�VF����(�.�sA M/-[T^4sVeU�3�UY�_P87�|Nǰ$��Ĕl`	��|qŬ��b״�ʊ�����|.��̒ҹ�G�K
�+�JK\�
AJ���B7�2�8�hn�� n���M�4��~v�3K
��\e�Ӌx|,*/�^)f���D�@wziIE������ȬB��ǿ�3A~	��p*K�+�PYXTQ���//��(�(/�\�X�i�~r���r�+���j�����b ��h\1�U���kn㺭���+��g��Z�	@�g6�p�>ф>òD��<\�q񐜥�_�>�݈F���Y�l����Τ��UX:�`�_�{��l�U}��/=X�ڇ�@�
��z,�h�o�3qy���R��[�P5���`�[|�͈T�k}�٘������	YX�N�`��-/�C�\+��\-�e!Ӊ�u'i!�d%�#m�EF/��}����\��1�E�aNiEm!>�!�$�E�	���'(.R��U<�p�����̴��V��zVס݄5>��#� �	�f̩�z�sa��z��`8
�0��P]�T_�3|���hų_�l�����	B	�=��=k�,��6�+�r���y�ck��k1?������X�"�����SOV��
��um�f�.�~>2#d� ς��RV|���	y�@��e������;k|����g�������>����z��.1�Rm\]�>?���pᔕ	x�Z�k��ĘO�k�إI�c��S+F}}�i�t/K��6��ͺ�h;�ŗ5h�Z����9��&�h��
i֡!���t�K+9DK���<���U����N���^he���&F���E�A��}8����ǟ\���|�~��f\�إ]�ُM���M�Z���
_��C�nK^`�.�h<�:P'<D�ΙF�JQ~� �԰m<�
�o7
ye�o��X�u:����^�% k����׹:P�_Ou�s��}�6H��)��h��vZC��M:���kĕ�%��0�+�isB��A��A	y��5�z�<a���*�A�~��e��9p�'�ѦM���s���|U��%h�蒪���A]Ӹ�yr����/"�K�}����OH�����
/�ag��׭�<��ÿQX_���G㸷�^O��0�<�	�y����E�W;�xĺ E5S.��n�ļN�[�v
�P��Mw�{�O�7���jh�G��j|=&�̗�ᘥ˽A����ޢ{ ���q �`Ok�f�fp����7@���>�*q1����+��`�M�6�v�řja��\�u{J��X�U8�s�6=����(Z����[*篷�:��]�ު��um}Ѩ����zʯ��W���j���{cv��-�g}9H��b �f�ѫq]�KL��Zf?8����c]��j�F���X�ǩY�P�S*�`��S��J��d��_��B>W��x��] �/F�/_�ָm�T|��K�Q�+����l�x�Os0����B��|�
�m{.z�q/�������㙷g��j����sw��s.�����u VEb� fs�T����|�.�8�Y�S�]҇��|�#�Ü���{�U~��5lK30��R(0�$�a4]|�"1�Dy����T���rz
�z��ѫaV�K����d�����_зs����%��_�U)d��A�Aݙ) ��ӣ���|��R��41ƹ��Y�7�<D*����8�b�|����R�6P:Wӎ�3}��S�bv��ڻ�Rq�z��\�W����^Ӊ��N4r��î��N���B��?�������K�D���>Y�
-��+�-�Y�B�}\�!�w�����q����}��oЎ���ߡ�
�=P�B��u+����p5�U����-�q�70r�f��Yih��E�}mh&�y�bn�y����bV��'4��Z�
�����?�f����F��o��ӵ\��/+�⇿/3���1];6���V��FY��b0,-��l���zn~]�|Bl�^ۥC���̄�׮����:�:U}���|�[����v����d����g�<��ޅ5�z��qhydp�y�2�]��{5��E����6�mW�>��ց��M'��i�/�\O��J^��j��F�V��[�	�� Y�Y���2Ѿ��ð�Ԗ�`Fq%��li #<~�n�5�>��oG��E�R�KEb���]dq7J_�ǈDOl$^��V��l#w��Ƀ�a��$���,9A^!o�����gr���\$*����iM��t���<�3h1-�Ut���h3]K7����� �M���q���qP��}��ў)�9j��L���ѿV�W���]#ڳ��+�w\1�Z�g]�Í���`G�B�'_�_}����=7��^����g�h�����B7����+��HB���,J"PoF-@��Z���hߓR�6�0�&�������Q��ލz?�?!cD� w\��?�;x��g*�}?p��V�6\��͢�-Ѿ���^!��iB�'	��6@���|�0B�#�h�b��_�ī��י�ŸU�u��9�Z,�sK�_]"��7H��bN��G��-.�����y���i���5�p�~/ǘ_��:F�߰��#na�$C��k���#t��?���]�'˲F�6s)Pj�u��P���{RjY�k��_$>�YvZ~���m�q��M����o�Ȱk����>��
endstream
endobj
38 0 obj
<<
/Filter /FlateDecode
/Length 412
>>
stream
H�\��n�0�_e��!"�$BJ�#��5�XR�� ���5+�����k�lۃ�FJ�m_y��3��k�5Ӊϝ�TP��cP�[_��g>ޯ#_��((�p����i�n�?Q�f��9��kst�x���iAeI�n��jx�.L���������y�*>���:}�ס��V��T,�SR�wOIl��R�vj���������j	��Z�!E��B�P;(���$�P(I���P0�9�K�'���,�*�(k(,-�H� �H� �P�^ncx���%�U��a[� ۪�Nc\-b\�ŸZƸZŸ:�i$��eE�b\��
�4�) �]E��(9
9J r�(@�V�6�< �o��S�N������Z�������z�3���C?L.��
0 ���;
endstream
endobj
43 0 obj
<<
/Filter /FlateDecode
/Length 15831
/Length1 36636
/Type /Stream
>>
stream
x��}|Tյ��g�s&ɜ<	!@C �@HBx?�$$�@HB�If�$3�$���H(Ҕ"���)�"�ǥ>��Zߢ�֪ U/E|�ZJ�3��sf2	���~���~����k����k�='�!�$[AA�l�s�"��$az^~�srU
!��o�^ZR��><���^2��2�tAأ��uԒ򌬍)wo&��E��5Mv��/z���lmͲۡ�G���6�ֺ뚮3q	!�h�p���& i�p��5������������z������7���Qz�����ojY��'~��	�}�jt��3ϧ#d�Aܟn��pGUj�~=ؚ�M��:~fo�m���m�#��t�׻=Nwќ��F6����=y��EN���D�~~�9������B*�֨���4�@�͎&���A)�#��I�s�H6���������QQF+?�m�qe�'�R:X-�L�%I�����"��'�Kk��Fl>����m�&��bB?�}$~�ԛW��'�3���"��3���%+I.]BG�������դ&r���#.���*�ET�[M��;�^r��⺟4�z��%��B��6�Z@����?d��=��!�_$גv�]�vH5z���j�-���s����Ǔɠy�~Ka|����)��}t�P�rR%r#i�b�@�(�o�Hc�s$C�A��R�5a�	D�����p��wA��[��P-d�C.�)��&c�k������3��Zp���aD��|�I(f�� N�bP���$C�������c��@ʃd�an#���i�Ɵ�@�K%�	���{�͟��wA#�H�̥&�S��vbr�&�X�)�fM�G/a���D������	n�1����(�, 7C/�	4Ê�⺙́������{)�f�@��4ĩ��ҾB�hK���2g�E6F��*�����Q��z|-1��i�U�-q�����@��� FM���	�0�Y�[h�IV�B���Xՙ�p�&7�m�F��lB�B���9d�V��,h?+�)P�x=���_`�8L%U��T�;	���2��${L=5B�����m��	X%w�9d&�^i"��y*�N+�4�|H=G>��f��+�JG�DS����u�t=�vE�(�h��@�ҙ��W�H;���/��p��{�ĈE4t��d#���_��#�-��{�����s�d���K�!��ڂ��Rh��9}e|�0؜|�s$�Iޠv�>���=鋄\��n�J*�
~��	��=B����W�O�*�(��4B����{a#wb>��	�����LWÚB��yX��X֏A3�!w4[�{�%�(;�V��׊>��X���A�I��U��Mܤ�$�CH�6��mq1F8˫����1������5���Ŝn5W�^߇�UX=��7$%��?�B.�0�Gn9���܀t[1b,�s�b@,Z߈rB�aW9��!��#�OŘ �\�#��v�VK`�vrzOB�b� i�j�E����o2%@g2yX���>�6��k8FZ���oHo���bo��O�?�s
�Å'9 V���Eo��c��;~����6D
�|�p�O�&����/;	!�і�t�X�n��/�b�}P6����4%�1�3D�A��%(w��h�����F��H�!�b�R-�`_�1�+ka�[�վcԁ�=Ԃ�ܟD�� ��~�M+h�A�j2����R&xt�Χ��^��|L%EH��-D�oF!���}� �����??���}�k�!S�s��r����GN��9]�z�6B[S1��A � _=B6c��A`�Z%�l���]���]��&�5"�j�>���d,�i9�V* ��_-q�e	�@P6� K;��v;��P�@C}g|���:�h�\=���C��s�7����������ā}�X㵼W��kB�lܕ�5�7��Z�x��M�� ��9�D�h`8�DK�5��	]&�,h*��nS���<0���B��٠Q�����t6�j*QӇT�I���+��NF���Y�J�F�H.�B���i&M"_�� PK /}Q>�=<$���c	�GU=Spdu+RDT�����kֈ���G,�RHA1�H|�r/ȓ����wES���&b�&�}���-<� 8���3A����햂e�Mxd���<�
NFDg�q= ��a��M���X_�/	>���G8?���Ew���Bg}�8�U^nF��G�G�:�:e}�>V!��F^Ōk��/uz:��J�2(���-D݉���)����~CGs�}�O��u��7\��Z���s^97/�A�H�z��+������xj�k�#d}QR�\���d�n����B_	���긞������?N�����BB:��G�h?� ?������ߡ/^����jd ����ЃX[���픟�&�m� �#Q��^@w�Gpf$���{p�K�݀�8�B�Ŋ(V��K��Q@!�&�3�wԧ⚄���)�}p̈́�����~O�g���� ����4¿�H�J���%P'��,��Ls���}_�g�(����:i p?\c�w聴;����ɤ0�.7���0��
�%OO!v���5=����Fk�Z �ۍ.O��}��A5z7��s��!�J��Tyk�aGY� W��Pc�"�Z�vU�z����%��(�a��)��	���wqz�B�΅�3�;�w��nws =[���{{��q�|0�ܟ��{�� +0S�['��*}�C�O���h}L��{�	U _+<Iq$�'��;U�����i8���?c��F�u�DE��݀�vq>s�U���3���0Q}gD9!'�T�Z~y~5��Y����-�lV�s�8�qPy��/�7�F�s�?���M? ��D�3,N%͈}�H��%��)�W)�c��7�\�����)���;CWຂ���{��� ś�!��z^��]3]�������.�F�^����t=���*��zI�*O��G�y��{Z����"6}��9i>��$�K�#H$��q�ޱ��.x�۰��S����3�n@��>�h���ň���x�D�ԡ�?Z�|���`W��uv k�����X�C��J��	����i|�g�M��l�٦�,#k	�[�����©ƃHl	l;����"���$�G����y$V~:�JG|7%�M�g�vDtCqJX�S/�U3!�p��l��_�	o9	|���*r5�v$�_
�d�lE�uX�����'BG����&������� �0��a�24ǁB&x��n �܍�c��!�$}�+gbg�©��I��G�	(!����9�O�mX��В�]v�Q�[�Z�L��߷ ����o}�?p^ji$v�r�q���� DJ��	�y�*>����x�V��p౰��a9�"]H+M%��h$����<�������������(r7�w������\H�X�r�W��i��U��8β1��|��(�N��}������ e#��c�
�Uî5�e����?��k����i^!�����<�,��������a���3��}�{�_i&�_� %:���p�Ǚ�!�?��}�%��]��׃�eO��������=�|������U�D�%���E�G|o�>\g�
AǼ�hO\C`\^�{����wҔ��U���|����-�5���ǌ��I'm�[=$��V�!�#���B�<��.N��h;_p����[8�ݐ��$��~�sr�~� � 1$�2�c��(��T�3�\ߞ%a�D�5>���&%XU����H�tae-��?}>�v�hS�6�hSc�iƺm|�\z���إ>��o<����q����6))��︌4��L\n���HH%f�1~9R�8����#�$'RR���i��LEB�Fⴚ��){���i���������'��}}���|H���t�Tȿ�Ig$Cki"��Nb���v�_�_�y-��gCCb�����?�X������_YTEf%i���Rr��`��*�K��L�qk����҃�+mG|��*��2���p�%�������#�f�V�>��gR�_����*d��Q��'����d�+\|�VSo�+����rNI�Hk�[�����SO�'/�_]`����~�=1��b���ǲأv��=r����Rv��ߋ=��}�W�]`�g{ڠ����g���W��Z+�y0E�3��ɖLa�u�@�՛ݿs�r���?�{3�'��y��s:�y��,e�R��,�]g�]`�.���lk�I2k�g��l��~��M:ksF)m���{b��q�Q�=�lC��6Q�;�ݥ�;�?�ܩ��w,R�?�֯��=Y�c�#[�=��vk�r[_vk$���ݬ�u��.��]�KY�`kz����j���� �7d�Uh�*���g+P�����l��Z��7�y�OW<:�>��Q�^�\��i�YgM�����Y�Z��!Yi\���K��,y�5d��Y=��;X.uV��j�3�9tV��j��W��:���^�,��5�lA�?2F�Ǫ��<�����,V���r�R�ʭ�lN�R���F)s�Xi+�Y�l�R��f;X��f�lfa/ef;+��f\`�/���,?�������b��YN�:�M�fWM�P��ٔ�VeJ�le�&�Q&������>l�Zy��MȖǏ�WƏg��ܸx6vL�2v3:V�Fǲ�Q�J���B��x����d汌x����D62-Z�F���C��JZ4K;"܍���d#��gq7\S�G��G���yr�,6,���R��+)CX2.ɳ��fH<˒b��,6�6F4��Pn���U�c��$�l ��b	���^J\������V��b����D*}�Y_��<9>�����@.����bǳ^4Q�u��d��,%��BmT���R"W��ET�p�	Od�5R��5���<Ģ)!�,Đ�	-�p	CeU	U�0��هd%�)G(��+��I�
Kf4h"#1�����#�����{�t4L�{�a����d!���5C��"����F�l��l��,���gP7Qz5�t$^[�$k��Xd����6����n5_ImҫR�ր����� �{�=���MF�4g�89F�(���I5{{�a��M������+��9A�&g�w��d�;�W�z*c#�Qc-�!��\ si�s�$���� G�Zi��X��qVZ(� m#'��t�H��x��m�s$9�����E�<ySlsC!�>6V�� �B�Vޑ��\��6��� �	�u�.5�fX�(g��Kp��iF"�z�\��F4j!��5�(Q���Z�IƱ�gF���g����=(:yP��z�txY��?�했��xT��T��}�3���aU �#�H�u��㯀ƹ)�deR���>��#4���4�'�U[}���q_��ݯ�:�s��u�+���<�z��@5�_TǙ,�ԩsgΝ�:�����:�F��Ƞ��>��tp��;6ftָ��Ăm��[��t*M�ܞW�V���w�2b�����+��!C�#9���C������I��
yBH4�ݛ�C�"E�ePx"�M�#g�'�3�d�H�1��R�A��TJ�ز�~'��Cv�~T߬��q���*��0��E���A&i��K � R�=�P�u��uѮ���O�D�����A��|�c��Џ����=13;f�4��ImL���R$���Et�<vP�E�R���X�����W[��c�j:r�����/޻g�O��hp���p��z��Fg�O����}��;���(��9�����ь��#Tq[TI�!aZ��cYǲ���Ν����l��{��qM�ߤ���1Z�2V�{t׀�B�5�D������2N��-Ȝ�C���;���;x���w�i����J��,'�%��pc��`ڲ�a��FV%cʩ�c(�̎��d�W��$�������%�I������B)]�]�_(�JWIW�\z��Vz��Hد-��H�6��2�x��'���mt-����;B׆n�?g[B��Mf�B��>J��<�oY4�`XE��8 �ŒZ;a��^���Aу��`=x.]�أ�Z��:��Rۅ��N�t�?+��.�-���f���	G6��ć�Id����B	��D�ͤ0��8�|)��0�꯯���S_�y3���4T��ޡw��?�Z��~��q��Z���^_���o�W����u�a.xJ��S�zK}b����Q�1Jx/���^(���pr�[�
w���<Æ��%C�B���30*n K�qܞ����ֵ��t����-��e~M�c�0�ޱqi"�+JJ�H!��1)C���*R���c��z�o]sh��7��G����ش��Hj�|z��>�H�?�V0�t�Q����9���1tTEY��i�����`~�U%���F2
�'i7�T��I����HoSI���R ����3�	r3����p��������?=j����k�����w��q�,�nmeT}��O�id�:��I��'�g�Ƥ~@S([�Py�O�ڶmk�ܒ;q�:����t��4���ɇ��=4q���c2v�(�@�e �"�X֯>"�>�q'ma}d'eE�YSk�@wU1��`l���Q�CqT���o����c����6}G�u�57_w]#{N*�Ǚ=�j:�����H��u��.$���NK�����Z��ػI���z���o�jJ�G���qjjw&�0CYg�>=uV���m}]{=����{��_Y���,�{����L��"�_�W����^��t�O�ǖ���n�
��������:Sn��7O��6�,��z��U�̧�#��������e��z��ɍd����)�GRS��8-+F������c�N���:eL�_��Z�Cc~i��e�W� }�;��,Zx��yh�_�/ZT������X��ɓG����Rn��~����/��~�?�����޸����Q��h�6c��E�G]GBI8��[i#�T�-�+3+�SH�%"���c�:��Uq��Q�e���΁���Iʣ�m�OЁ4Y����c݉�&���5��[l/�$g�($�������k�'���}Yl���@=6n2�SR
�E��T\V}Z?��a�6[|⟿����{]{Y�����h�F�Z}��	�Ag˗w��5�a�=z��{*�'g��/.�F�<�}��wI��L���j�xS�y��E�o���ݺ0��g��&��wr����ԋ}vo�r��QF��I��+V4,Y��s���Y�W����g�'|�I��]4�^���x�^E(�\�bͤf�FĲ�0��!.���F��勡��6�a�4H�>��u�ݝ�K�#M���)�1lDZZ�Ԕ���y��=C�s(y0��pM��L	�,a��C��0k�@���;ve|}4������K��o!S��E����&�����9�!��a�(Y�=�Flt�����jM�R�S#�ze�f�N�KMH���:0�6lА��A�.s�ķup�V�!��qP�h�#UՎw�;��)��&�o��[2�9{��>~��W�Ș�'�f�ؔ_l��/�d��)'LI�Iٵ~ס�Ѝ�1J���D�D�F��&����E�D��u�e�S0C��6m,��/=F���
+O|��~����':���9q���|�NŘ�s�����!;YE�"+XUɈ��F6QU�M�Q,�{�QTƩ,S�<B
1����T!�1�R�:3&k�R�*��j��P�ߟ�����O��4�˯���܉�Ζ�ׄ�{,��-<j�xC�ɽ��$�"z�J�<�i/���X���i�:w���\���fؽ��t��5�M��7����9_>�~�I:�I�+Ĥ ���p9�A�^��%�4=-���Kz���,�ճgٳr
`����c�$`��*����W�
\�+p���W�
\�+p���W�
\��/`����'�F���:��+J�pg�%"��g�w�\�+D#-f^%��Z3����^3o%�n3z/y��G�1���Cqw4l����fM5�	��2���Ay��[�ͼJR�~:!$��#3o%������^)Z3AꭏOs�Wz��[l�jRmY���m�+m�-���ޔf+l�I��46��x+����uz�9�ay�%�����z{s��k�{���f��������p5���m���^�lW�˖�jt�uz��f[V���F^ϫG�j�O��õ�������ʗ��{]��g��S�Lov�d,oXڐ���p�Hw׻3�j��^g���y�r��:��jg�kyj��H�����m���F^���k��c��hk���&�g��UۓJXX������E�z�ǉ��<���#�V������4[��fo^isc>��U����0J��-[��D�kj\Mn4�Z�A��дmX�PIR*�9lv��U�`�x�`Mk��������mh���q�����U۲:OJ�x�n���Z�d�����)x��!�T�����,oh�w�����s ��c�d[�h��I�59��b~��iAc��13\�׉y@��j��ch�Ⱥ��[LՉ��׻�.������ӌ����e��l���%Κ^b�&��q5;��Iaa��W��9��	F��j�4x�R>+�.0�l�z;��v�Z0r{79]Ͱ����q^Rl[�J��֎�����6�Wr�M.GCm74{cL�;BrCu|}�=૵��9�ކ�f�F]�Jw��w�j�/�����s$�����Az1��y��W���:D�8�{,E[��re��/'��i���qxmI������Wؒ��Mj���	�`5q���.�2WC�1�������W7:y�!?(���z{����Egsw�`�.w�Z�"�����$C��ͬn+[L�(���{�C��f���a-�����7�nC�i�Egc-gjF������V^RP1/�,�VXn+-+�[���gK�)�}R�m^aŌ��
Z��W̷��r���f���J����m%e��٥E��(+,�VT�WX<ݖ�~�%���م ZQ"���
��9���e�f�6'����b~�������, �[iNYE�ʢ�2[ieYiIy>h�lqaqAFɟ�!@hZI�����3*�Щ�i�������9e��8�%��&���Kа����g��r+�+��sf�\;ӋKfsU��T��r�!JNnQ��D�V�S8;͖�3;gz~y� ��)N�:x�����e9Ei����i�<=��O�-�{h�H�;���<N%
��?&dF����4����r:%eV����r�
�9e%`��'zp+�O>y�&�|�x��ցV��)`^~N�s6.j��_Q�t�p�6���+5�g��Z�	���7c�e"{��;���ߒ�L�������~˜��^�J�>\ܙ,o����m��e�{^{#C�@+�K{#�ylv_P���i@�垆8�����U�V�1����Qz��qz�ة�9W�����g���fDaM��B}5-��>��V'�; 8b�t[�F\�Wi u����#5$�,�	�\5Z�H.ڴ/��8����PZH��>��m�,@�+:��v�e�Cn	(�%�hQ��vP�-m�s�6Piv�ג5�w�ۄ��'�rA�S��V�H�g�:Ђs�E?���>F���(���{���>N��7�k15��m����7f�eh��v.\=��)�z����Š-h�\-E�R�+P�M7ʊ��N�����ד�.�^����s���}9�������t���K�lh܎\0��[�xȿ
|���}���m��.f�Ihu)�\����KV*�5	j]�kЮuNS�:1J��G��S+j��ь6l/M��6��ns}#�@�Ŝ�a�,5���4[�W��j���M�~
���{c7�法d%Ib��b-�W�U�>vS>�k`�M�J����V�����a�F����߂�`�9�K'����(���.nB�ak�e�-��?�w��f��p�*�:Y.l�^x�S3M�,X"?}O7�4�m:L��o�����E��#- g��R6A�X�S��g��R�5gp�XtK��h��G���j��m6%t�����&���U�NH�hlǍ����P��!8n09�$Vg�ً�P�%<C���.\�	��KE�����ֿVܗ���lBf�9S���5C�'�_f>]bG��s�$����l�6+���p���4u��\'+�7��� ֲߣq�[L�g����K���<������W+��E?�D�)��� mԉ��]���C��z����S?��)��9�Y�]�ѥ8�<'��멗K�f�{���p��1=�S��ԍ����L��鹋8M��6˅T�?��bR@�=x{���dm��)��T�u�
��\��X�چKh��d-�^�[��.f���<�ϗ_1������k�����bHw)�k[�(2X_I��W���Ὼf�f�l3%�:���Dc �=�St�^
\gΘ�/�|�������n���5�bM���qJH1��8%�� �O��:�7���h��w>��Q���j��<�X"~H�f�(�磄Ӷ�{~7�A���'Ub�|�8޲LО��"\��v��_%�y~:�Ѩ1^�x�M��-x18�@yרݹ*#�9���2Пa��v����O���� �&�9BG�2�9�;^Z�k�x�V��G��m��� ��,��c&���Z��y�¦
���l�&$����|�Y���Ĝe�n����&^���.?�M�_��
179��뷝���U
�r�J����k��(в,hV�	}�y�牑r�F�/)��Z�ٹ�u�G�.���*�ˡ�|�/��X(d�f�֠iؽaEAڝ&d�3;��6�#t�]
c�p���0f ��ӂt�5����N�u�����2O��|�*G�uy@b��69��0�<V��Y଻~����������3�'���<���k��|�k5�c�k��u߹��Ǯ�48�L#]�680��tѶ�G��R�?{Vי'8�����?%1}W��>�m����_��ӍX��J����L��ڮ=�86���=�א���ѓ�_�E��G�^B��ۡz��b�7FY.�-fd��k5���U=NŞ����,ߧ��o71�TB�<�L7�z��|֥�㻰���e}��$�3�:���aθ�3�x�#>���/�\�M�	!��g�	2��=��$L��Pi��S�Iې�O��;��o�� L^/����ȿ)������ȟ��$��������=�!����W�$���|�0r��&j^AQI�{��$�f���L��8���F��F6�[��4YH��`�$�Wa����
�QF�.�Kd	),�m#cf	\$��"�b���ϓ1��9%]t�cM�O��ӛ�6-�-��2�"$S�oڙ�g�JbI��C��]�����ڌ��zX�6����е�}�.!�eh���7���}�N"���JK:��>���=T^|
I�DkΩ��-�8V��:�o�oÕ�k��-�]�"���9���%"_��G0��<J!$2��L`G�����cl��M������|�k��T���(���1t�ݹ6P�ۋ�1�U����(Tz��{�H��7�렣�$禮�GK�k�����W�$�������H��I1R��(��K��8i��+͐��
i��X��%��B�I�U�K�$�Kۥ]�^�tHzJzV���������tJ:-}%}+u0�����1Kai,�M`SY��J�\��U�z��Z�*����6��l+��v�}� ;̞aϳ��k�8{�}�>eg�7�<�eY���89AN�����y��-�Er�\%_+;�%�[^�U}3��Fy��M�)��ˏ�G��1�e��w�����Y��|A��#_Sb�x%Q�W2�q�%W��+�e�R�4*e�r�r�r��IiW�+����������-�=�C�rZ�J�V�P%5D�Pc�~�MMQ��,u�:U�Sg���\u�Z�֫�j��J]�ޮnP7�[��nu�zP=�>�>�����W�W?V?UϨߨ�U�"[�,Q�8K�%�2̒nc�dɶX�,e�*˵�e��mYf�s���p#_CR�^\/lu�k������|+xJ',Prt���M�� 8��k�"=�T��z���<]���ǒ��W\僧��}���#�5��(�@���|^�����|<L�X��(7pE�g��Q�;���L'|8=������
�l��Jc}39_�1z��n��r�������;��v�a'�1���:���t^����(1J�����XP.��}�|�E��
<O�Tl�#�,Q��cz܇Y�[|���D�\��Ǿ	��6ʫn�3Hwt���v����s�����M�21k���A�u�����$�����dK�.������|��i�C������ȗڣ����cz�+��,�Cb.J�]��	|�X�:_~�����d�\�� ��������~�R`�^��Z�B}��:,�>�k��� �u��ho�/��߄�	,�� Gs�.��}w_��Q^�[�,F��]sI�f痗��w"�+�E�T�����@y���o>��|kx_�]���q��;z�����*�|TPy����|;��@��{�;�����eg	�ߋ��b]����#��G��E�� �K���N�x5�E��O�z׿��x��)����D�O�+ݩs������?m	m��z�����&�莥��B΃^����� <C8/���S�zy���9.�D�,����������L}��
n��a�<yB�kD��!���FFk����R�4�զhS�rmb�ڟ�3�S��%9��������F6�U�b��Q�f��QRc�УdzȀ%)��K�"�P��E�v�|�|�|bu�׼�����������������7��r�e�[�Gz�z��m��|7����Y�Y���0�t���_�oi�$I!R�+��lR��&eI��R�4S*��J�j�^j�Z�U�Z�vi��Y�*�vK����a��y�%�5�������tF�F:/�Lfa,�ű�Ć�t6�Mb٬��2VŮe����2v#���g����d{�~�;�c�e�{�}�N���Yv�]���ʚ#�ˉ�y��)���ȹ��X��ȋ�Z�Q��+`9��wɛ�vy��K�+��O��ʿ�_�ߒߓ?�Oɧ��o�ERB�%V�ؔ%M�R&(S�<e�R��U*�J�Ҭ�(������e��U١�V�)���3���K�k�q�}�c�S��r^�UYS��85AMR����u����Ej�Z�^�:�%�[]�ިެ�W7�[�m�Nu��_}L=�U��/�o���'��ճ�9���XT�f���[-C,�-��q�)�\�K��²���Rki�x,+,7Yn��e�di��������#�R��y^�f)����\V���������2x��4���}���O�nE�g��*��HY� zT� ��0]%sϖ����R)��J/`��G�f���]CRU^�)�+MUyD4��ҷ���2e-c|���� >-��'c��r�4A�{���Yz��AXZ�����=^AHp,E��s�c�|_f�</�&p��A��'	�+�b���y4U$sy��p���;�J>��
�ӮQ�I�B�-�e��*8�H����
Wp�c����W�WXxT���ڔ3�!
�b���G�)�.�C�<�Ű�е2���8?�]�
��*84���G�R^.�H�7rE���� �y�\"��1�{�\��B��|���$�
�8rA��cZ� '�)O��s[B���Z?Ƹ]�[Yp�T��
��6���4��;-:LT��D(�ar�ۉ4^��ZR��ת���qac�B?aWù\R:����
�����BI��w���hNA�R`��}��x�$�Gz��3=���V�̭w��0p����kb-��,�;�8y������ȭn�Xw�`��(2�.��'��Z�Og�>|�	����1`�2;���*�bG�oR��a���NWy��Gk�s{���)fv��cU�:��2�_(���&������o�U��C{T��)�O���n���(�+�	��ƹ�O)��t+�[1}O�p.�G�Wx�Q�\%f�x�Vqr[R�:-��@I��#��
��S�P�h9Z�	������*?���Z��)3n!���P�W��y�ZA$/�<�-��G�|z�7�Ÿ��
�tXP� ��:���x��L�{@x�G��T�S���瞍>�r�xX�g@��K�b9v:g�s��<�D
V3������j����T���VjWk�d���8�&G�q�7�Q���2�ǈ2n":�i��q� ��t:�N�ٴ��2ZE������2z#��������{�~�=B��c�e�}�~���w:���~'�x����!�6��\\{1��\����c��ǃ�uA��6��
.�!��_����	���	֌()�!���� �u?\�����:	��.G�U�B���<�|����� w'���鲛
�sD~�9֬�x�)~�j���<2'�b�H���zx�����w�Ɛ��򗁓q���dͥ�d�Ag���M�&�B?�������2��o$�^�H��32��3�q���!�̅����dI	��m!Nv?�E�,,H����F�X6[������I�u�u/qY�Y&n�/��$�A��k=d}��Z߱�K�[�d=AV�_�OW�x�Cz�H�B�j�zb���-�UHk�nG��St3���H����"Fz�y���^�7m���89����&����{z�H�=��u���*�w;d��v@�}��0dyr�F������Sr;����c��X,�L��M����K���w��@�-�v���j�Cʿ+<���K�>.�*�nI����(A\D�;|�f�w�� ���MS��w2�`�?��S�H����4680�8�3���1-���1K<k,��ĳ�j�1�a��F�|�gO��?sT.�t��2�uZN���旗O�)O ���*��J<��O ���j��J<��
<���J�������I&8���چf;�khnh!3Q`'����F2W��MNG����������,�qĳEN]����L`��3�v3�k�x��g߸�o\����8����X�8��T�ǵ�+���'�aD���O������nĩS�l-W��
��Z�V��is�ڵZ�V��kK�F�Y�h˴U�M�����]�Fm�֮m�vh��=�>m�v�z����S�i�ֳZ��jZ���Yu����цkI����U�։���WD˃�/�/ ���j3�b�B��j�5���Z�ڍ�Z�Vm��AۤmѶj۵��nm�6L;h��~n=c=o�JӴ-J�Ո��ٴ��	�"
&����8#Kr8��o�H��
|ā��$^~��i�1]���k�k��ͥy�������n�M�W��v��s��!m�����ֿZ?����w뗚U�h�Z/�O�Ԓ���$������H�L�;b�$��]x�j�)�D�X�	��i�gk�O�5�D�c���J?a��P�w���	p���B�4´��o�_0RC�Y�V��+W�z�_�~>5ʸ�F���D�
endstream
endobj
46 0 obj
<<
/Filter /FlateDecode
/Length 317
>>
stream
H�\�Mj�0��2�t�ؑ܀1��/�C���Ʃ����,|��z&�⛙7Oh����hOɻښ=u�(��pu-ә/��6%�[�P��}c)	�z=���*
J>Br�n��Ag~���)v�\h�u��Wk�g�iCeI���襱�MϔDٺR!��������2����1ţmZv��0��J*Na��F�˧��ܵߍ��SY��.�[��v���ڃN ��`��=3�z�P)9*evo$��G� �,2����{[��؂�A�(h�/��{w��9�Z�2^�r_��s�M��:G��<m��~�`gU�~ ���c
endstream
endobj
47 0 obj
<<
/Filter /FlateDecode
/Length 10019
>>
stream
H��W]��}�_�ρ������lC���rYB�&��C.���J*y$�K�mu^b3j����q}=��/�������o������������')z���_���wJt��ןO����	����z���R9!-|���O?������"��7���.�?�z%�8^z7�A�=}�R[�����oR*XK���O�SE?�j���WW)-<�������;�w�k@�e��}~���3�l��>������3>�k��1>~�?b;�}��.rĝ}{�,����b��(���/
�?�4
��h�r1L�h������R��Nj�^�"�/���:����� ߩ�������٣�y%��g�W��G���EH��i�7:���iV�N꘹ӏ�"n��n�P���v���b���_��fd"��RF)����Z������ �~�a�D� �&�麥7;^4�c��W4¬����n{���ê>~ ��L�S1n����(*\� )m��"�
����̈́��Eu����ԥ�-٨�F���T��\��*�19��y����lۄX�b>fj��C�n1uMǽ0�d/�ҼٽOqg"�0 $m�+6�����_.��6��6�+Ek]rÏ}?�ӛ7��M�#���1Wf�L�����g�pϦj�/6Δ�g��Wv���l"ڬ?�,�X��Ӵ�!ز�8����I��Wj���~��jw-Ml0\�����K���BL�~*W�U�˲�_)�鴿RbݵM����⻊/(���0��X��@$@gj�n�tjM�P�� 7�O�4<���4v5�7zVy8��NZ+a�������!{6����du�٬�Ǖu��+6�ޛ��M�C<��;����a��s�5���ަ~\�rSO�Zo���M=��pSo�V6K�զΑPV	�����z�V˦�g��,�{��˗^���OXx?���c�i�J"l�+����A��ٛ���7��i�>����;#��w�@�����Xڋ��覛������\W���	���5��y��+�����ߗ��-TcfY�O,�2�e2�W �	���L��t�R��{�HWڋm���{�Z�_��p0�T������$�e����Pa���!M]�6���]�|�H�[���/���8}#���r!P���o)&-4m.��[�hc��?S��g�|=�����f-���R������=�js���'��Y�f}�R�s<��{�D���f�o|��Y�~Q���:!�p ش/��$z%���m	�N	2���1F��%���ϕaM$b�"��I�mKI#�.<�*�y���PrZ�`>��Y�@�b&�0�:����lh(;����
W*�潹��(�A�и3��,FI��[Ɇ��hiC8�-��Ɉ�A�M���+9
~�'�	|? ��%ST��u�ԡ�c�Q|K��y�ʴP%?��� ��AM����q�r�]�M�0ٱ�p���?��(5ٽJl�Ra��py������ur&�5�nv�T�T�X�ˍ%�:=5�xp~������W��U�n�|������-T�(B_��<j&�����຦7^1�X���Kd�T�Z��QƟ��{��'R�����?��V�`+�1��9����E�6�Q�-���y���Ny�R��w_!sª����۸�R���he�n�8�^��Z'�����w��ۮIY�֮@t�X�R-0�%���E�\��Uq�YL����Ju�0���Na�B�f���<��sݼ2�	wcu���}�E�:M�l�g�Bs��	Zn>�1�;�>��q�-[���u�zl�Q9�,���D�|h�1�l���BX�s�R5��x$P]*��Z�R-4�Ka�Y!�\�O�=Ο��VZ)Ne���F����W\������:����N�V,�w�=v��3j�C��6�[NN~�|���{-F���?f��A��z�� ���Á�;G��q�u���'�#�Fw���Q��o5:{��Qx��V˯�g����۾�8�)��<h*��S�1	�MI�7��GoO"�V*1Qj�[�<~93/!B�>�YGSP����k��ܙ� ¯L�.�5�����U��?͎�(�ͤfʀw�i�Y7�iRu���8�yc?9��R�'{���7Nq�<�-}����|�+�C�E�=i~�[<8�N����]���ʮp<�C�ð�lW�Zt��]��7�8��Vz�8��{'7�V
8����n5�Pp0�Kvhρ`�t��7C⸃����`��B$ƾ x�TڗO��w�@�b��.�{ȼb]B��>�Υ7�;-��xȹtA�/9�~�g�	|? �u.ST9���1����%�E�z�н̬�Se�������;�	�R�hm� ؔD����i���V����Y��$�fV�PM^�W~�`��pT����)�p����B�5��d�Q�+�:��Ԯp���3�hW�̦��o��`:�O� �ve*�*���0�p�<�j�]�jѹ�;�i�T��)]�0,ͽә`+��~Y�j�W
�)��M�Ϊ5� [�DtV�F�"��ŨH��tb�
��	�e/t�5�*(���v��B��zŮP��N�v�I�֭0��̊U��*ÚWa�wp(��'nK\֣�ܯ�(g��/�6;�� �mnP��;� ����%�e�{G5�։7���n7�(��!;4g@�UL�z��q�d��ū���@�OA�:����H3�BqR��P���xş� iU݉1�Z��?1AʸfP�-�H'�	� `֨LEP�T8��h�#�6[��m�B���_����������w6G�:��ʹ&a�Ms�Nr4��.e��&�6�b�j�8�B�U�yc�RifV|�T��[%�"��
��GѮ�A�!iiW8�CvE��hW�kv�����t�� f��TUv��a��y��f��բs3wbӾ�����Nȁ��w:l�V�/Z��J6%Q�)䬚���J���H40*!O�-FE�|m�cT�N0-{|�g�̫P�L�GەN
�B��Ba�:)��aa��+�!��@���]�xp0��'��Y�2A�]�x8+�P�a�ٮd��ns�rOo�q"�u��0q�1��Nn��pEA��<jJ��` ��О���0�o��q#�������H�}A�J��/%�J3�B�2��]��6�yź�(Y}���.��s��8;�޽�\nk΅���u�� ��GT9���1����%�E�z�н̬�Se�������;�l�f��4&`3�Bަ5D��!Z��q�B�$�fV�PM^�W<~�`��pT����+�p����B�5�����Q�+v�¶t+�!�2@�O^ť^����jɎǁW��,��W��N�O������0 ?iR) !���zF�,��t0�7Y�~�sM�ƽq���־$�P,l�g�E^�N(��~�G\딚n4:5-$ɣ��tB�u:�2jC�	%5G��Qe*��Ma@&)te�'�L�L�kD$�/�L�2�y�$e�V��CI�� �LRvioI��Gf
�T(��n��.�Яx���7��d:y^Q<�xx��|�jw>����w��{|>����2��ц]`�.Q1��P[
Ln�Zr�xV�ós$�G��C_Q{���#D"���2�*�T���Q������ ��$��Kw?��s��=M.��f������%�O���� �L.�K J.7�n�#�v'��.�6�x��ee���ʜ��{�IX�f5�&Q`[L\)�f4��*ԡF����Rw�h_XIt�LT^��2�r����+�K���a%m�<2P�;��~p�q�ͤ@�o�n��� ��p���&`��?oכ�(�\�5��]�55�v8SsQ�e��Q���7!覉ѝ�>E�|��亸�Q�1Q[k��m�O�J�/R�d�''Y���
�����y�*z�,sΧU��2�3d kɷ ��7���uJ�Yõ���i���=�LZ�!��g�
���Dȇ�ݎ5�M�Snd�-�՚����7�O���t���;��E��L(�[mG���T���>�{��շ�����o�f� ���ͦ�?_�7��b�J����m
p��!����1�k!��l(�Ϙ��C��v��zM'��*��j��������Ý���5Z����/�+p�id�����K�yZ������-�B���Ջ�S@��^��WQ�l�+�,����\_�ؖ����L�=?#d�'[�ဟEF�����vS`{��}���s��f�ͻz���p��*=�V�)��0�l�]y�N\�+��~U�U|�Tf��rV$2lG�$��҃�m�\20}���&����N�oR?�T�*�dXa��X3�|
0s>L�u�Õɨ�Ӂ`f.(�+<�0)=��z�9O��;�A����pH��ө�v��`�t�&���X��X�T�K�����b���x
.s:3y:V/*�7�
+<�S�K��
O��%�S���C�uF��Ra����ˑǥ)��4��{�w��
�	��xQ>hQ�ap!�8�ܱ��AD��Y�㙣r3�j��6id���F�g�_��ac���0�2��~2�e��?�/ 2*�y����b޴�(zj/�D^S�ߎ+�P5lL;���^^�8���i��F��'�`~�>��ì:^��*�����6*�8�����/}�� �[?�Å�˴�V���d���b�F�Rmy)��7���9��/�q-� �Z�m�zz`���i� vP��Ë�]�h$	�1��2M�4�J���:����>i��2�ZeX�V�S����,�j���*�K���WS\)��m��-JY���\���X��FG�A088!����!�4�v�i'rȊ9�J�͚��h�趈�B{�]q����OL�Ș��AW��jFi_^�7���T��~��ܲ׎\w\�>����T�i��2���ث����ៜy;�82B����tj�ZO��
՚��a<�ے�_4��>�D�*_�Lb�f�I�BN������C�hX���`�u6�+��`�+	�wدFCO�&L9���
��Kz�2�.7mii�W&�vV�gA��^�9)��dx%R��G4�ɍ}c��7��}c�����/���EEqZv�q�kO&����c.��� m����k�y�>JOm^����A��Q��
U���1Q�;|�,�JN� wҸn��8�=V������_FʷD嘪�Q��!-vpȰ��^R+wi?�TX�Zn�̜�ṭ3�hi�S�l�Wŕi}����۸�@.de)�h���v6��-���7)k6��_�ߑC���?�?������U���?���L݌|�i^�a��r�P:rݩ$�X��c}V�	��ZnUݞs�rf���K2��v¹�p|��p~�EAMCT�X�Z�V1�'Q`[��&��ǓȰB%��9�ؑs��u���ֹ
�����Ծ�oy���I�ʻ\�F&��[<3�v��T��p�����P�q�^�J�5��!n�j�}�ҲUw1i^P��Bc����$�0�xH�1:��ȧ,�Q�b�k��ƾ�o��ƾ�o��������8�;m��*��'��/�S���ʦ�35s���g��t�
+T��28{$���(��0�7¸����aXK�ߚ�7(M���3���Sae��iV�P-���"�v�����s��L���V3 ���R&˄?�f�!�?wo"�^�m¿���m��}�yw5�������|_�b�n��%`]I�%c_�x��#��zsA�_�|������}�v�၃�7y[�����-��j++�_��bgs{T�iT�V<���}�퇐�F(�1͘�Z��R�`<Z�3���#3~0���Ǭ�ZS^2D�%�%=�"o ���:��c�_���w� �o��
Gn�8����LEV�EG\+�I?�i��:*��
���W�����օ׆G�	wHio��_T��-�$/4���?���>��^J�T\/\h�O|��Kd[��z_|u��Hif"������A{�S�@�7=��X������.��	�,:�a<��7ԋ�F��覣�@���z�Y���i��	�!K"*:�'�L5��!&ӓ��	�h��c��'Q`eJx�����=���&9���\+�L1�E��Z��Fy%�Q�;��U�w�ӌ�
Z�A�	+Ҫ�P;��_9�h�#�����yQ��p!~��jD�G�We�m{�<�o�uq�C���b��9vX��:� &u���R�-Q����V�ìU4	U��i!'Q`��z����BVN*����^I���K�!I��$���w�"�&�zK	����9����[��k��H��;(���s" ���7O���U�m^���9��h�F�z6������S�)��+��ܶ@l[ <˸�������a�O���ŮS(��ESH��)dT�
�U��@�X����~�����U)�׆���d+c��*n�e�o����4v��OzñdQQ;��M����*���J5aU�3)�=M�WNA7�%]��IЯ(�g����7����B8\��K��g�4��ɽ�wW�Tt6l���(,R�+V��R�J8��?��\Ҩ���9�x��M��i��;3�E��	���k{��7�xc�T�3�ٗ���a��!7̴:�1������[M�ࠗ�M�쬕���:N�c�V��;7m�	�j[���/���m�γ�^�">��N�,k�Y�	M��LH�P��N������p�i%����'��;i_yN�.��y=�K��eON*�g��U�?����p���ŏw[ZC7tC7tC?Aׁ�u�ٗw\`�Bֹ� 2z��|y�\w�l�~11�3��j׹ėeg͢3�w5,��Ȥv|:i��N�tM��Fئ^��$�g�����sW(�i2�*f���ς"�'y&�����
?�;P�om����	��̖���p�L7�<�p��h\?u*M���TY0.4��p�L���]���u&�������H^�@��ڛ�_x�q���v����I�ˀ7��D@|�V�c���4��#>>� �@OUp�RA����������5Upk��
QSA2z�U�+WKe�Ei��+��E&��T��tNUPJ26�\L������D�0�dlL�*H�QSA��+�,��aB0݈褐r2H����K*H�:����~�
�5����
�s�k��J��c<����rꗡFn�Fn�F����%�ǔ�f}����>�X-��ʙ�D^�$*2���'�Yu2��'�L=��ܔ=�T"T
SA��塨��r\H��6�~��K��{���
BE�$��By���������ֿzC�^��H��HY�	淦�q�*��*@O����؂�מ�n�n��4���K��+D���詖>�\-�eM{P�T�ԅ�=)Zu:��'%)�z.&�ܔ?�d"UL�4��j�#��	�vd�f�TM�0!�n��$P9�ʂټ��%$y	E�xo��[��[)��� {�*��T�M =U��+d�_�����ZS�f/QA�5$��Z�r�TP�]�6�A�Ri\dRO�*X�Ω

CIƦ��I47UP;�H�����ZI0j*�b��%cS?L��=TN��`65�yII^<�ó��T��&��RVA�eTUA�X��a��t�'��
��/D�������[��� W��
��S��\�Z*(�.J���^�4.���
֧s���P����`�M�N&R��$ccj�VA��
jG�Xaf�����F|O��A�,�M͸`^RA���
���u*��D@|�V�*hDM�U*h<��S�W*�T�5tC7tC7��
n�^��\!j*HFO�
r�j��,�(mڃz�Ҹ�
.�*X�Ω

CIƦ��I47UP;�H�����ZI0j*�b��%cS?L��=TN��`65�yII^OU�h}Wu��oM��o���Ɔ��4AX%���S�ƕ�+�~j�Fn�Fn�*�K�]�}Lj֗ϙj�c��r>QnQΔ'�
%Q�����dN}OH�2�L���rS��S�PY(���+�6�<5�S������i"�u���馂PQ(�r1��dxyV�	���]�K���)�]o`Xh�G�<�X���	p7a�_{����Z�����D��B�����j���U�>av�ИR����~���c� �<�9�r(o�I��/���}g
�����4<�'N�[T��)b��L��s�vU �S튛$�&�Xab�����aB�ny�����:�4���F��R�|�"W�0�{2�p�"�$Vt:�[�[>v:�X�ts�S��.��-h�p����^�����'��a���LY'�q�seXUB���HO�����/�ޗ��+�v�����qŨ��k�g�_�q�W��Zv?ˮ<���F�)����� �tJ�i��"���%�w�W4p� >N��9���-�[���'�Kyk�đ�UX=A"^�C�����@5���K�\�~l>BFt7W
�g���F�V���G�ϕ4��jDC��&$��ժ��A^�hx����U�~�z:헫i��ʾ���+��������ί����Tnj�8�q9��1�7R^u�,�㐨�G��̎�+��.h*S�|c٭�+R.պO����毫-]��Ȕ|{?w�;

+/�τ�k楫�|�E�w��l��F{���,�|�~g��T����7�5�Ub~G��E��Os~qĪ���N�ϫ)�4�pׄ�x�o�n��	�Π�v��W�[��C�����~��i�:�#��W�<�m k�p �lp�N�;�f@�觝����ߵR���x� I��rĪ�$�\��s~O��=�b�i�~|\ܸ^��\,q���p�sq������	�RR�;a�3/����3_o��"_��d����x�E ��l��'ol�	?o�}|{��Q�E�,-�O��~��hp_yNcq#5}7Ϫ�#�l�!�@?�t�j�q�-n T?��i���[���h컼ϔ�a�L
�>����#�>��!���21/�ȗ[�KD�0��
}!�z0�]g�=���+3���C���_��6�����@���d��d͢��HA��b=���	Ko�C'X�����w;���rR(b�i��f
��B0��~�G�磁���ßF�Xa4S���L��)�6��F��CKB,i�?�`�e���"+{;:e�<��	K�N�n:���V��K���YF�K���4KiI�ݲp��#�*��u���KXaZ�'^8ˈ%E���A�Я!Re9��gJ��rAM�"���M�y^��&�lR�����c����\�x���> S�ʯ���%�)��]�a�{h%&(�w7)3��fJp6�u�X?]�islӉ�u��#�l�sU�|�`[���J���y�pQf0���n�ˡ���O�A�haB���R^�.	������Y6a��V~�(Y�am�ΆփPQ$`M�a~��'h~�Ȫ?��������B1
7��PQJ�=�#��� 6�TBW�S��ډD�(�$��C*@,wp�J���z�	�ڻ` �m.O%��w�*�ddf�Ó�l���p�ٗ�ܨ19i��)J�[��I*@�k��2i=E]P�� T�؄���O���PQJ���������C���>A%�߇6�2�/������z���w�S�v�LtI��f������%~�T�ޑN�۸��{<���-�A�'�Za�C�m��~���J�Ͼ>|f>�s�3�����j����&��Xc
��nT��"ucq��鵇z�Jb	�7|�y��X���n�%�G�)�.U:- MK�G�~�/U~�Ŋ��X�����@�Vf���ds
�[I�$�a�Ҥ�ۦ��IM)����_�W� ��
endstream
endobj
51 0 obj
<<
/Length 960
/Subtype /XML
/Type /Metadata
>>
stream
<?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 5.6-c015 84.159810, 2016/09/10-02:41:30        ">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:xmp="http://ns.adobe.com/xap/1.0/"
            xmlns:pdf="http://ns.adobe.com/pdf/1.3/"
            xmlns:dc="http://purl.org/dc/elements/1.1/">
         <xmp:CreateDate>2021-12-27T09:02:53+05:30</xmp:CreateDate>
         <xmp:ModifyDate>2021-12-27T09:02:53+05:30</xmp:ModifyDate>
         <pdf:Producer>Microsoft: Print To PDF</pdf:Producer>
         <dc:creator>
            <rdf:Seq>
               <rdf:li>Acer</rdf:li>
            </rdf:Seq>
         </dc:creator>
         <dc:title>
            <rdf:Alt>
               <rdf:li xml:lang="x-default"/>
            </rdf:Alt>
         </dc:title>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
<?xpacket end="r"?>
endstream
endobj
5 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 6 0 R
/C0_1 14 0 R
/C2_0 23 0 R
/C2_1 31 0 R
/C2_2 39 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents 47 0 R
/StructParents 0
/Parent 2 0 R
>>
endobj
57 0 obj
<<
/Filter /FlateDecode
/Length 16631
>>
stream
H��M�����gmp]�Z�`fl$H���E�d1g��OJ�ӧ�ԥ�v�r'��~��J�RI��_�����~���?~:����ç������Ɂs����[�~y��y�τ����뿦���� ���yJ�Ӌ�L~�r�������O�N���I;����N_�N�<�	=�9��ӗ_'<q�xbA�2�/��o�a�#.�\��/�>��"�z��<���q�H{}�_�����k3�~�����+z�5:��Qƕ?�֬b���^�ŏc7g/��_C����g��Zd�|�F���q�C9�n�������`��`�i<�t�n:��F
����޼�m��F�*rk �w���)Z]�]Q�R`nE0�����k-���!"�T��I~�o%Էb(�����8~��oS^oG'V�ϥ}�7��=뷖���<e���i�@O(�D!Ӻ��=�6R*�)0��S�9�#�e%�k'�2�=ˁ�9�t�<���*�'/`0Y�f��b�����m��+ s*e��3�� �G�V��a����1�(G��P�Q�~�P�|�P *�x!�"x�-�q��%3 �S=\�YXeatf��.�,����Qx�k��S�]�4*+9H4-��*KX��m$c�,�Q���v���U��\V�s
��}x�f��H,�ph�	G	�m��c�%�&�t`a��A3J�k���jI�_e����?���H��:h����2�|�^9&KL�8X�tP������U�_e�s���?�=J�<,�<J�ͯ�J�
��Ű����*Kv���X��ь��얮O�_e����?�=Ye)q�ph�����q�%�&k,�U:hF���x�J�*w�u.���0�+%�ޱ���<���HC�L�8��q�0���y��h�_�vH����爋��h;�F�(Ў�R��U���\���q���Ջ�3����};��I�٘,��Z�ca�rG3J���z6&K�.��Y��s���	GqZ��d�c��c������)��v`��?�bퟅ����.�A/٭�`4bj̎�1��(��#8��dy1Y�p����l�ﺆ�F��Z��d����?c���Q�d�H�Ie��?����Sȧ�ë��0ۣ$��m���N���U��\�ן�1���F�S��"U��L���\��;[ k�� �ml���� �x*�ծ{c �G5��o@�J��|T 5C�4u$���� p�p9�
�#x*���P�� 7C�"�datF�F�5������5��"���/����o�=$2�]>���1�d����J�(��	�<���*K�.��Y�/b�ӊ���]t4D���E�YeIg@͚c��3��2]6��S�rݧ���j�����z��i<��@�$�6V�v\隣��M�r!��y����H�PD��G��Q&�����֔�Ƣ�&]�}P`2]�d��L�<LsgV�Nϓ��F[6�$�2�x��@�^�P�S�ė�ZKsy�u�\��'>�_X�h��v\�$,�m,�\�I-ǔ\0�u.���2��˅���:���Q���!��Gӛ@0Ghc�|\��W���qDw��A:#]R�[#w\�ZwT�^wT�-�9.�]����e��"`-��*!�.���!`:�:B3�pfC ދ�)<�.W�Tw�R��� Ѽ0v��.p0��<�U¨N�@N0�[�0]�Y	D�)����UX��"%���' % ��: L@��S���J	�)�J���� ��k,̆�w"%��*�?O�ː�֖� 2 e��1J	�)���
L�NGd�	�0�c%Ƀ#�c%�����蔈^���Ŏ��Ukz,�U��N�@v׆P`� 0 cM��ٞ2����]@T�H�>�Ȫ P�@X��P��:C%��U�K:sk��L�����Sp��7�R��� �5f�G>�!�;m�O�V�;�1&��m
�)�yVJG�钀NƜ@7��;g�8I�}��W�S)���n��ހ�5=�*T�D {��� 0 cM���9�n���vs\@����0V)�:=O+̑���\d�	�0����S"z>���;zL�FT���0F��;%sG��I\d�	�0[��%�S"���=	]��&��X��D�l䮁� 0 ���Sȧ�ë�0�c%�"�:m
�����2�9��]�u��)����.	�d��;[k�m�����E;K� �T�]������)��
�/�q����x܍�\�&��"���H8.��i2��!Э� 7G������r9�k��=k����ݽ/�?~~�D5N@��D�}N0] ����X����s�OsG������+~��͉(r"�J�^C��#m�<w�J��\ b� ����)����3��N���){�:�z�ٴ?��q�~M�}�@j�z��N�r!D�y���B�{��Q&j_�+�ʳ���R"z�w�������Ukz<LOog�Nϓ��V��Ì����5f�?�{��M{pդl��pss=�6�L:��/��I "����_6	����2��d���G1��馸\�9�s�|uQ���8"?~�	s\?,�0�k�l>.�蠴���@��е��i���]j���x�-��kAuKcz\*����p��%3�UB=\:��C�tnu�f�3�.,̆@�MSx�]�l�"�¥b!\�A�ya�p1]�`4n1y��Q���`n��`� 0 ���Sȧ�ë�0(S�Q���	��� �uJ�0V)�:%�Bi׷�`� 0 cM����N���W%T��ivR���r \@����0F)�;%!];[A���鈌1f{�$ypdy���_�.z*%��w���tAo@՚c�?�S"�ݵ!�.�X`a�����ȯ�ݸu��y����d]7҃�i2�=T:c���&q��bN`����\R�!��R)�������X��Z)��Z��  q)�˘li�ZR|9�~�D���Z�dei�s����.��{���X�L�X �M
�R���~V�  q)�˘��6�l;i�_߆m�z���v�øЛ�Z�A��Q+e���ƅ�D�Z �|�>�� թ�9��	�5��j	���%�FK��&ƅ�D�Z ��K���z���1zG�����1��RX9>�aK¸��X@����c�^)Ġ\�^D\Ld� �U���@rT��2\`1.&2�@�%��m�Ǉ �~[���J�@���&>
lq!0���Hct8�+�^rh�{�,���eX�-���j<A�ħ+���$%R�Ű�����r�z�3��4j������*<މ�]���������p^��)�r��^*�H�W41���h��ar�e?o	li��C��G����� �Z8��@��Ϗ=q2���4V-�V�%���e����h��S�g�I�D�?�r��<��2 ո�� �� ��|e�@�����#���K	N��5S��x�8��k��=���|r���]b�q�0�!�]�ú}���h�Xe�>�_�ů)�ǧCߔq�m�����7�	q�	��JLL3b�j���%�ɣ6�� ƅ�D�Z ӌ������W�ʜ�N�:ă�sLߵǷ׈�;��� ����~� ,�o0�VoT����u9�gg䀸�ޣ#�N��[�C,�>uOKr}-_�K��z29-A�ܩׂ�)�~�;/��J 纳4~��uZ�B͟z-.Q���y'^1��R� z�-���h�w&H ��HO���[��R%�Kea��(�O��\F�+&תa�JY�dZ���[\
Ld6��K�����	�pw^6�?�� 5��5 [\�L��[�k�j�,��~|˃��k�N 8���*�~�,�P.��q	2������^)ļ�l����d�p��m%ˍ��m%���zHOUb������-.�&��z0\��Q+e������R`"c- ���2�rIq�@��;��?�d�K�	�5ת%�JY�-�B߽�->�2��p�ZR��UB-�z�\U���-q	2��������#z�]���$)��E�3c�Ѥ�+e�X�WQ� ��]�\��/�q�g��I���6l��S�X/e�6q�7Q�փ�Z��Z)���� .&2�0ܯ�g���:�6q	2����Z��Z���|�%q���R`"c- ���]��B��b���P����p��G���D�Deؒ .&2�0ܽ��c�^)Ġ\�^0.&2�0\�P+e��xN5\`!.&2�@�%��m�Ǉ`��m%P+��R��(�ƥ�Dƺ`�F�s���%�F�S�a@|�eX�-�6^�i�h9SK��ғ�H��fwG{8���j��Δ�GШq�����*|����%�iJ>/�_(�n	�%�r^C3#�Ke���Q��!�E�3�p��o�O�[�p��C��G����� �Z8��@���[\�L��A`�V-�E~gu�@ɴ��i�������|�}Od�)m"��! .��t/� T���h�K��=_�"0\����;�W���V�q�vˋx��96ϗm=��;�a�!D��>�ۇ�Om�*~��k�>���z|��׎=���������Z����U�~3ø��X`�]�����-t�k>�ղ2���ɍ���;�_��w��� ����~� ,l�%����;��`��1r>)�˂�X7�G�(F �g'����!�D���y	�B��d�y	���ץtb�J%�S�p�9+j�JP��VvZ��O�O��j��kޯ�J���n���R� z�-ı�����	@��@z���K�r�*�C\*seG�����q�5a4�bb��Q+e��>H����&�|ɱ|���!H��a|=�� 5��U��de��ƪ%�JY�5��������� ��	'Z"[%�¯������A0.@&P� �ƨ%�JY ��f+ ���d�0�~[�r�(r[���В�+�^�T��+/".�&��z�ƪ�JY���B( .&2��f��<�%�Q� �B��� [\�L��A �UK���@[��U�K]�\`K�֒��!���%:O���CK`\�L��A �~��>"�W��zO�[+��`�I�W��R��j .ts�6���a�b'M��۰�~@OUb����ƅ�D�Z�X��Z)����0.&2���k�Y�p�N��a\�L��A �UK��^/�7Zw�0)0.&2���XRt%��^�aЃ8*�T��0�Q�蕲����[ƅ�D�Z ��K�JY �Z�"�B`"c- i�z@�����9�p�Ÿ��lɗ˷��4�m%P+��R��(�Ņ�Dƺ ���\��zɡ��Tm���|�%��XM�G#ș�t傶����D
�6�;���@�WCow�|<�F�����P���N���4%���/_���O������R� F*���p�q,uF���-��@xK`K�?��?��o�@��$��~~�	��	�5��j	�(�;���  .�=o͊O���D=��&��=O��@5��KA\ �{��E �Q��P�Å�_/%8�R�G��m�����-��0\���ɹ�:�9��q��ð�������C��D��*�Y��,~MA>>���s�\b�<D��󕘘f�<��j��K��G��e)�q!0���4�@�\��n��_����9}��u�g?ʽ�k0��%`2�=���7��d��mP��J~0���2r��%80�u�{ԏb�yv"�ߚ�`I������W/�G��� ��drZ�J%�S�9SJ�6w^8֝� �ug%h�T��?-A��O��������Fz���_/���8��~�Z7Є�MI��i������Oj*9a&�.��C�3�D1A�z3�ı�����O	@��@~���,o��J��).��������y₸�Z0_11�Uè��@�c`�� ą�B�!�}-��8��)Hs�?EK�v
D-�AZ"?��4�@\�,��[�X��Z)�Nm|*� ą�B�Z ��-��j��Kt�J}��"������^)����V@+]�`��R��Q屒�뷧�]��r�:�]?�A\�-T�� �U����@u����X�X@��)�Kn)��Z� i�'7�<�dei�ZB��z���~�T!.ts�G��m)���Z������盟Z�dei��ȿg�J�@�ߓ��#���d�0��K�W���8�Z� .ts�������$����t�~BOUb�\��ƅ�B�Z�X��Z)Ԡ��0.2���Ϝ�z�Ҝz�ø Y@Y�@��P+�^��3w��R`\,d� �����+�^��: �I⨴R5��4F��W�1��Ou:�0.2���(pj,�+e��k݋����� ����RȎ��T��B`!�Ⱦ�T��� �9+销Z�h��8�g�G\,d�{ ��z��K	�<���[�q)�˰�_��<V��w#(�^������Da�����Z ǻ���)�A���[ܗ�W�<W�}_��2�4��K�����O������R� %���i8�8���Q���|/~!~'�Hs�?��~�xD-�Ar��U��' .@P� �ƪ%�JY����5NkHsl�*Z"�Lϧ|T�i��_���g�f�i�:ćJ�d'n��KN�㼚4&:�q|����ex�;h�1�?��B���e�?Dz���e�6����f�GT�X���M"� .���z�f�;��j��K�a���Y�q!����4����-1����r���%�._n�wOy�a:��1��;�X���J;.�[��YZ�-�v2�����F�!��Vp`���?��9�|�,�1�`{ݗ Erc'��dGm�Kyc�F|Fl��L�+5��@a��x/�����ߖ�R�[�x�ڕ�Gi\1#�Ke���f'�c�+���ɟ�4��$.M�Y�r�*�S\*sG�����q��`4�bb��Q+e��ȏ�L� ą�B�!�}-��8��)Hs�I����a�9Ձ}z�����Y�Yw������%�J��]�P �B`!c- i��	�6�p��V��8��2�4F-�W�9�oyB �B`!c- i��s$�M#�O���S�X���Q�A\�-T�� �U����@m�q�T1.2���x���[�;�� ���w��	�dei�ZB��z���=	@\,d��Lsl�sj��Kr�*�~z)0.2�= i����+�^J����U0���d��o���5�~��
��|]�a7!��1�k���w%H������G�h�M�7!ȅ
o�~����b�%���4j��&͑�Qژ��>mK�3�������TƩ��7!����K�)�t���r�4�D��M1�L��úS�Ƌq��Q��}��<���^���sM�t�[ 7��M1�N}<|���{�M	��4���M��H��Hؗ x
��`wS�Ke����	�M�RW4L0d�{���;�G���w��������	�pɁ
���{�dei�ZB�����M��I �B`!c- i�-QEK�� �������>-��K�@\�,ܬ} �Q��P)�~�<��z����B<�r�ڼ�sD��o�~.��ypn\���e�?g^��!���e����h��d������� ?>��Mg\6z�0yI�|�%��9�̘'�Z��z	<x���) q)����4������l�iW,g�zQ����]�8�1�p/�pX,�{~T;.�[���Y|�-�vPu9�|u_��z�Ʊn|����`��ȗ���A3�y��}	R$7��/Av��d[�F|Fl���b�%��nW��v%�����ߖ�R�[��e�c1��x�4"�Ke���f'�c�+���ɟ�4��$.M�Y�r����S\*sG�����q��`4�bb��Q+�^��T��؎놁4ǆ	�%�l�g�NM|���X�`�h��3e��[�0!�h+d�v�4F�W�����?m�kHsN4L8����Nn�|sK@\�,��A �UK���@m�m�M�����#�A ���i���i;�����z���w��I�Bo�j�i��G��zI�S�:��?kHs���΀��~'%�#�����A0�QK蕲@j4γ�&�K]�\��������+�^.�Ћq��P�փ4V��V�%Q���I �B`!c- i���P+e�(�`:V0.2��ƪ�JY�9�4	@\,d�ג����4�c%�P+�gxą�Bƺ �Q��[ЋR��R�S�x���/�s��_������-��G�,��o��Yu�)}��s����Y�����q����(F "�,rng�v1�痱�}	R$7�=q_�쨍�yc�T��z/(��a[��hl=�K�~��^��z�� �� XЬ�$J ����A)�������؇?�tl�����x�il:D��r��y9N�iRD��$:$O߶S\*sw�YrA\p-��n�nz�,P�q��I �B`!c���<F�̷#h���݄�7��ʯ�����g���C�>�w�S��Վ����a�#@��n����]lM>u����X7>G�Q���s����-b&?�޺/A����÷%Ȏ�ȟ7&hT��z/(�r懷}	j����/A���n/PǛ�r$�8���[)�$~T�E�F2�lhT+�ŨV�ڕ�c�}Ǻ�9��F����_�oA �ڮ0��J �ڶ�QmW�v%�QmWլ�R���2��pY`\,h�9)�DS�B �F ����_7ˍ�:@�~���%��˶+y�������$�JhLM����n�8�(p�Ҷ"N �ҵ�:�c�3(e�F�%�JI S���8��h`�^��! �2�_�K\"qEg�	�qA�qM��0�RÈ��@N�;�a �&2�����č5L�K>���`l{��8�i�`�+%�ZMi�~S�8��h`�^ :�!u	D,�~�[�/��J�贄\)	��<�0�c�3e�fh	��]��G�_˒��Dz1<�JL�Lo����i��G��~	�59��`�	Ld�0��?�o)�)�럶�e\���f�^�#�Y���i'�R(;}' q. ˨����W�=o�8ݎƝ���~ٙi�A��� jG��1y@��(��X��}4�s�gmL��e%�N�+0�J3Ue=�F��JI #]��q&0���4�ʰ-N TU�����J�(��X)	�,KgmL��m["|5,����r��-��`r��8�0jsa���+%�@clk�n�8V:�Q`i����-q��g�0�'�z��Eg5��AgzUm=L��?b�$P�8Nc�	Ld�0��?7�!�S���p�,�U�)�.�;.�3�	�6�Qj��&P��N��3���� ��좀T����l"��W�\@�Q�4:=`]6>=�+'��]��b�O�'��I�/,���{X�s���/K��c\z.b�7�q2���4�bg��6���;�#�&2��f�aE�&�U�O_A���;]|�m0��7s�ki[,�"0��E����=��C�,~_��*��Ly!�J�je���X7�G|(J ,O/���W�hlm����|V؞OKp| �J@C����%�������g$�q��OG2��J{ �MI,��Q1� ��E�;�Z�ʾ�ɨV^�J�1�#����ETE^1�1�����NKp�j�%x�j�%8F����i	�QM�@,�~q>۾>�@�Lh��$L3�?lP�� i��k(��h٥�+�2a�`j��aq�6CV��4J�$WJi3�:���tĹ�DF[ Ҍs�k�-���7�b5��=�3�A&P� �F�%�J�o���}�r�w�����f�axK��a���|���2�`�h���4����8C�!+cb����Kb�$�ÿ�7�\`"sD�S�o�?�4���Bɕ�@H�I�q.0���H3����2�}���{u�/td�,�4�x?���EX�He\ƿ��g�Y����)+$��ɚs�&h�c�x�h͕��y�p�;|4m������-Ɵ� nϏ�i	�+�S�)�ۗ��9����KP�qaS��R������� �&4�sK�D>�����Q����'G�WleC���<&M��Bg�ʶ,�Nwɕ�@*&��vgmL3��ܶ"N 9���d��i�ZB��~�tO_�� ƙ�DF[ ����r��C�0�_�L�0�5�����a�f�ʘ,��N�%��&P��>��8�L`"sD�S�o�?�4���JI ���� �d��4C�/�}_�i��:��Y��x������`�9�--�ғHe\ƿ��gY|��7e��ϫ�6��Ǻ�>�C�3!� ��Y�W�hl;n��o��?���m_�y	��{yV��L������`�VP�y	�3.l�{�X���5!�g�9	�1��^���Ǩ��%�4�j\n��sqd�1*sa���+%�Lm�@� �du�#�8Y��p��X8�Dg�	߁@��L��A �VK���@���@�	Ld� � xK��C��_��ט�eZ����e��?�0bb�aN��1!��N��R��D:�n��8V:�9��)��`�q��Kb�$�y���G�L`"���f��쾯�Դ_@�
��'��dj�-��6~�iK��֚T�E`�{��|&���ڛ��G����3�}>#C����Ekr�<���Ǉ_Aࣱm��%�l�����q۷����v� %���y	r0m+���6ս@,��>۾>�;�@�Lh��$���{1��`���O�]ڵà�F�!���#w�G���a�贓\)	�ͤ�X� ę�DF[ �s�k�-���7�b5��=�g (mL��b���i�\@�Q�4��["�����p�;L�K;��F��O"�{�0�h3deL�fh����\)	xk3b���8�������Ǐ0Ͱì��X)	��<)0�3���v`��n앱�+ 5�P��BG!�����~�m0��a�5��������L mw�7e����d�8f4ın���P��J�3��~��>�6�|^����Θ��q{~,NKPLv۩���Ll�)�%�������g5����Ņ`j+)w�>�3�	��i��g�P�a�;*~�ӟ���v.��6:�4}gq4��+�b��+%���� �&2��f�y��m	D,�@r2������d�i�ZB��~��O%r�3���� ��-��7���+�a2�\�ad4���<���qD�!+cb����Kb�M���}*k/pę�D��6����?~$ i�&�	H��@ϩ�	@��2�= i��_p��R�~u�/T��d���}�m0���a�5��������L0K��ܛ���^��l��8֍��֘�yz������Gc�q+�� x��#�?/A�Li��	��{yV��Ll�r^�L�
j8/AqƵ�+�b���sք0`�Lh��$�����
?f>F-�d��U�˭;{�#�,3Fe.�F�a�JI S�;�;�sYF] ���k	�-���Ht�q����J�(��X)	�jJ۲S' q&0���4�@�-n|�G�pe���/�v�~�[6)�3
#&��Y��t]�+%M�Q��X�c�3�C ڜB~��� K3�0eI@���5�9��(c�	Ld�{��z��?��+ 5�P��B�!���=���_.ɍ�:�{�ߏ�oW��h��&m	 ��4�;Hq�����u�O�����R� �7��|&$Y|C'�lJ>�lx�;33�|�nr��P��#�w ����#��Y��/�����a�+�h���qc�3[ς� F|ʾr�6
j�Aq�Z2��@,�A����O���K�&h�}Mw Э{1�e��e���ϲ��Kˠa� ��G�`^:�6����t��I�	$)4��K�&d�	�tG���ƙ% b�H���lm��9�	(m $]��+=��.�;2uW���-|����|�d~L+0eh�y��J�~�A�AV�I���D@�	x���f����D�Sȿ�?�� Iw�0u��X)���K�&d�{��;����2�mHM����� �L����^C���-%a��T�$���$4�	�>��gS�)��dG|�4�i���h�J�'��r�3����E<��c�}Ds~,�EP ;��,H	"��Z�E��QPþ����,K=n.����-}Dg&h�}��ܻ��nU|�۟�G�%3D������[�S�3��lY��+E�@h�ێ ��	m4�`�y�8�D,���	���	(m 4�RK��7�<x��	P����&@�������ϐp�&�cZ�)CC��§a�>`T��f��a�0C;ݗ��6L�T֞��32�Sȿ�?�� 3L���H�"�N�����h� 3� ��۷ 5=���5�ӽ���=��*��n)	k-�2&A��%��LHW�I����diN���j�Ӻ�=�CѲ�$�@��]�G �Z.5� x0m���"�J�7FP���R���ײ/�����EP���g�X�qs�B#�34�>����׽��mT\�%ci�*�ܺ��u���2.F�a�J�@P�;�;D�d2��0��~g-���p|��BtdJ	��b�H�V(md�� ��	m$�@ �>C�*��ט�qiQ��7o2��e�)L�3���0I����+�J����P�KuZ��E �I!���4�8a���"o��we�32�=@Ì=���ݷ 5=���K��0=�'�z�O�����R������|&4Jx&�lJ>�l~�;33�LtZ7�G|(ZΑ�鉼�>�>B{7k�A�`�װ�A4PZ��1�ٙ�gAJ1�Z�E��QPþ���,K�eП���)Dg&h�}��ֽ�2X�2X��g�ц�eP��01���#w0�N�� k/�4�N;ɕ"�d a�ھ���L�h�a���ƙ% b�H���lm���	(m 4�RK���m�꜀LF� 	3L���'�?��'L�ǴS��0���ҽ_T��f��a�0C;ݗ��"o�epDg&d.����"@��D@�	�tn
� ��	��a�x�Wƾ� ��y u7\���	U3�ur�O����R������|&$J�Ϥ�Mɧ�-�:k�c栉N���E�W�8�ח���Ghf��}�]��E����A���ֳ %��Ѷ� hwװ/����2�9�R��CgX[I�[���L�(�$f �w�/�ݪ�η?Ǐ��
+le��6:�t��cKt�p�\�-��]r�H ����32�H�ц��qf	�X8�	��[����6F�%�J��w<~�J���L�h a�Hy���gH��	��1����!Lo�����2Lfl���R$�i��32�hs
����? a�	�Gg���G X��A2 Dg@&��[��[����
���R�qÅB�?�����*��*�o)	k-�2&A��%��Lh��L�٣�1���n�c毉N���E�u�8=��W���G�m���"LK�� �sZo��@vf�Y��ivE�u�\j�A�d�Q�b���9!���L�(�$�'#��
�3�Qa����B#�[w��.�b�aT����4�\)j{rG�蜀LF� 	38�w��,G ���>�; Dg@&����0J-!V�j���#@tF`BF� ��%����;�5f~LK0Eh�͛)Ya
����6Lfh��
�R$�<x�@%v�N+���D�Sȿ�?�� 3L���ёG ��iӽ��P���Rn	fh������q�pG��W��ur�O׶���R������|&$J�Ϥ�=ʇZ;�f�����ߋ�N���E�H�8�׷���Gh�k�A�`����A4P�\�#(���z�1~��z�6
j�AAٌ�Ƴ�⩍C��@,��9g!��Pls#:C0A3��v��f 
�Ѳ�7䥍W���`��X՞ϥS3n�/	��!r�H����CG�蜀LF�Ch��@��C"��د!��)���*-�"[���8[�3����E����������9�32�#���z�~�
����-o2�����86B�/q������̏n?bEDO�<~�� �0�����R� �7��|4Jx&����������D�<uV7�G~(Z��鉼�$�>Bs�5� x0�s<o� (-~�A���ֳ %�xy-�"�Xw�a_ŁFu����j"��p�+�t�`�F�I�ؚ섀�f0J�%�d�������I�Kg��@)aatZB�	$	���-q����6�'�w���~-��v$�Fˎ6/��5�6��=�S�0'��a�0J�$V�J �\�\zG@&�N������)-G x��_ȥs P�@h��+=n>��'� :'0!#}w_B@���L���@������*�骰4�h�H��$0����\:{ ��gk�0:�)Wz܂��S3� �9�	m4�0�xg��
����~���(e ,�NKȕ"�`�6��}��ɨ��C�|?͟�4Cd,W��6���:u�k�Q��0b�H �����q�� ~7��A�>-w��M��]�m�?)2�Q9�5��4b$�����B@�q�4�!��f�CT��:B��n�>�ƩC�J���j�2v. q.`�x`�f�]����t��k��,�nq�b1:s�4>�WJ%�N��U
��B@�q�4R �s�۔��@>u-�&�h�s����8u�Z)	lE��1�oL�7݁|:��h)�8�!�}7oL��!j����s��R����� ��v	�R�7�rq!�˸@�P+=��bH����q.`�x`)��]&7�K�:�;�>{��{�>�8s�ܜ}X��+%���NK���ǅ�.�. i�˔�Z)	��^`!�oL��j�$�z(�E�$Ĺ�!C�]	0�0L>n����0q��`��B�*7q�B�ݟ�-�i�ZD��X6*�҇$Z�\����4R��q��7�2å�W����bt�bi|&&z]ڦVv� �tK�+�xJ��?R�8>�=e�5b�a=�mч�5<����Zם��w�6�.j�B��A �@(oH3�Lv�Z鱤��t+b��80d�O;�3<��j�S�N'��=|T��=j�=������s⑧&�q�9_ؚ�Ʃ5�JI���QQ�81�oH3�V�3��l�~��J��%�=�@(oH��j�ǒ�C���\@�q��[b�;̅�0�<�Ć󼞮Dz4oU��v��c�,Ug=L��?z�$����uH�3C�[ �|������Ձ|JS�!�3����xu�Z)	l=�s��:ƙ�!�- i>�c���Op�,��[X��Ŕ�q�e0zsA��Q+=��P~��0�oH3��[�[
n8o3\:q���70�,�3�qj�R(=��ޅ ę�!�- i���;�Om�؏q�c�y�@�Q+%�V�9�L����4���.�VJ[
9��J���L����4^=@�����y�5! q& ��]	`���m"��L�S@*ı�5�WA�3 λE �S�蕒@��u�X�%�,�iF�ˌ�ޔ�>�-�j�c<���w|�o?���������%�"��E�����K]����7�$1Q�5��N���0�a��程���H������ ��o{]��Ú�M�JP������	h�O�K���Z����l%�[�^^����·���xs�#�+����W>%a����5�a�����Q��ח��jo|T��dx ın|�sq�)!� R:���0�6�:�>pL0�{��n���i��}K��X���w�� ƹ�.��!�f��;��i���ƿ���u��=�n���?>_�x��ˤ/-S[C�Q��1��a-�s�b�F�+=��r�4�t!�q&`�x@�A@t�lT��e���C��7�m*3�:)Q�~���̂q$����ӌ��?e�/~�#��*a$1E`����5�`�����Q���K��TS�lp��0�1N���e0�������˷�? L@�n
endstream
endobj
55 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources 56 0 R
/Contents 57 0 R
/StructParents 1
/Parent 2 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [5 0 R 55 0 R]
/Count 2
>>
endobj
60 0 obj
<<
/Count 1
/First 53 0 R
/Last 53 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/StructTreeRoot 3 0 R
/Outlines 60 0 R
>>
endobj
59 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227150656Z)
>>
endobj
18 0 obj
<<
/Type /ObjStm
/N 31
/First 242
/Filter /FlateDecode
/Length 3970
>>
stream
x�ŚmoUG����W�oM!�z�jEH$4��
�d�+p�mb���\�ο���:�1	�g��O�:���Z���Жu	c)c	uI�-�,5w��ޣ.Q��U_��ʻ/��]�z��Ĵ�X�%ť���~�4&ﱤ�wֻ�]Ғ����k�[�k�K�z������]xkmc�#�ES�����(q]��QJ]�2T��5���aє�i���C8�ꫣ���:�_�_�Z�=9�_�?qt���������˽�g�?�U��ݛ7��?�Ų=x�߾�wX�~t�͓G���E�X�����ͷ��W?�Z����l{?�������Wo�������/������U���c���O:��<=�8��X�]].�\^�}�}=�O�d�Y���ӟ����/���7_�N�s����g�\�&�W����c�_�ݟ����۪5>9��>�����v|����鿖����hڳ���7�˫���޶�s���קo�4��� ���j�'�\B��x�=X�nM8����^��ӄ�7vt���[�]YAtP��WO���%W�vٵ���%F����/!,���R��Oi�;��>A���z>λ" ҁw��Z���`Z�F�&�{^�x�[}W|U��[K����}nAx�H',������m�#2���]D]�Ye��4���a�ˌ/B�&�h�ܵ��ĳ�me�,��-5��=�� ��;5G���Q����j�8�fA�G�>A��\4�.k`�h��y�J�f�T����hƀ^S�$Y�Y�%�%ʞ�^�"ۀ:eD��0�Z� m`74~�nRD#Ւ�C�̘��sGY�<�d��R�4��4�6 hj]fNh��A���;������M]8���JЇ]�Z�PƊiC�_1X�����$�`���([P����N��IF�$���T�K�P�eo �s48$��	j!!D�W)&B��U+�E@�#K;�(Z�d�F=��(#���;6>�!D-��9�嗺Z�U�)#y������s����}�X�\�J�#�	o� ]� �j�$�� "Nn��N_MA���":��L5��M��yӾ��\�.���<q����JM}eTd(ƍ�tx$!�����%��6�h�r^���t�ީ��$x\�x�֕�D�}���8׌�r��p	/͠����<���� "�x\x�����W�'&KBe��p!u\���>R	)�7��<�����f�(C��ZW����=`���oF�.��A ��+B�R;F-�c�q(�]n�k	��u.�#d��Q^�2Rs�;�C��pAsfO�/�ޝA&nF�Ê��-R��ULI"W6)�9��̩����yڇ,K��E�/��I�"go�-��2{J�����_�,�uOӶ���-Ξ2�YQլ/�=���Z6�[�/A�=�ԗ�18��!�P Ac;/Y�̫��E_��~Q"ۉ��a�%�Vğ���o��Au��V�U"��L���?��,iZ�Z�.�"nT�TL����uG	����.bGK�&S�K&PG�4�w���&4�9Ҟw�;��m:F�yL'm<s�T��1� LT�X^l��g/�۰>�c�}l��ā ae!�h:���*�.�vb�N-^P�n����Ub�#�a��@ʖ="& �<�8��"���0L����j�*Mژ��0��B���i��'R%�*=���L#� E��@Hm0�C%;��}W���fw��1�+OwP��y�GUFkg#5V�C���j �1j�uۀZHp��(����TA^0�>rԕ-���8�������X����n����B�;O��wĀ_R�0@*#B��c�!+�`uV����߬ѢiRcۂr�&n��7��⥓�����m�8';�³8橤zڳŉ����g-��Zb�fj�Էu5�����񩖕�HP�3�mخ�i��(��j5l�O���0k	m���K'	��T�I{�H�t�OO�J<:�A;�*+פ�6�%|hx
i�4E�Є"�Y���酉"����4�v�E[-0X�D�=̘��&=��Lb�y�p>褋 �z m.|m����%�Nod�Z������v��iBl`P)a�\Ͱ--)mc0�u�R&+��ՒL����^���蟩�����w��~�j�-y�.��N���bE��Zx��J��̧�p=J�%ñ�C��z�!��y+�4���]��vÇ
y&w��
5y��_�pV�Ôj[�l+F9�"w�P,�\vD�Q�=��C{�ѻ��ԭ����c�k��ʉT��N�.% HLB^զ�w�b�7���D2 �s5h���d�l�3�'�;lڊ���w��'aY#I�p��b4���T`�dիr�B�6]�
��$��Bt�������9*Um�$*�x�F�^�!�P�m������U�3̪��@>�����u�@R���LZö� V��2R�?w�DU*[Kq-�<��)/}q�ߚU���+�Q ��h]�e
�
�u|�d�$�i�sL'�$ǡo&�6B��&�����4�1IL��?����T�S�����o13p�G�B��U㓤�(͇X!�e/��}Ŋ;6�> a���]�;����8]�ǫ;8���0�I�F�8��
��$܌5��'A���hy�Uz��JsH�a�1ݰ7���,h��7L!RB�.����RB�P�΀d�#2H�*�޲D+M�\��Aov���gh9�ns�)ӗF}�^N_HLC>�H,'�i�U�[��R�O�V)��,�9�
�3��T��q^ʄ�
|����3Սf
o8�	^�
,+\`R�),"*
�s�I�4� ����o�U~���!P��$��\ Y#dk�$G J��i�̀�-fgaZ�	Ez�u�Н������*�Z1�
c�b�H���J����@�e}��\ �ҟ~�A�+i�l��H.+eK�|��\ �
dV�6^r�Y[Dȧ�Sh�@��>|��P�Npj�K�[�	H��`��K7¸P�|h�xȉkpR�X.�;�����f�ɒI�!AN4C:�2���9�g�(� 2##�tG�C�@��u,���)Ni��DaJE��+�f,T���7��mćm�L�3�<��ܰ���z����ʆj'ʜ3Hn3�oDP���ٷ��{lo[��$ꄳ��:��w'�z	0/G�N/4|˵����r��򌫙�뫙���8��>���ϋs5�k��ߍ{ ��ƽ��m��>�~L�Y���ɑ
G;I�5���v���ǥ��0J�7d6�<.5�8�%��R� v�8h�%?.q�3K�wm��o�(U߷Qj<.ͻ7J÷o��+�K(����x\�<.qx5K����Y��k���ĩ�,,N���Y�a�u�S�9[�~(?��<.qP;K~\"o����RY��8G���ln�,��92y���q	g=K��%�Y"�����5+���J��]O}�8�仏7��R�KJ����2��+��'���_�<zz��=~u�v�S,���r�ז��]ז���w�&�ؼuysgw^*
��h{�^���u�o_��y7����7i�\��N�q�q��&�]χ���&�����m��s�̄/����̟���q�7�&qS�E\Y�q[��|���|���#�M�s7��qe:�0q��}����ރ�.���O��G��>��7���[P�����x�9}��#P��s@9���Wd���;�(1�{�r���s�?=(�~tz�/��9�1��:�Xҗk�SZ��vO/�~����w��\�������^�Iɇ������c�yq~���zp�����_/_\J/�~X�{~�����6[v뉛>;��d��V��g��k����B��M�9r�}҈�RN<��Vs�^��6���+Uכ���a�oazw��\����pzvz8U���~1%���c�F�._��4L����o�
endstream
endobj
61 0 obj
<<
/Type /ObjStm
/N 2
/First 9
/Filter /FlateDecode
/Length 102
>>
stream
x�3Q0P0V06㲱���+�-V�6P�6� 
�**D�B��\vv`5!��
��%E��%!E��A��%\��@�F`�\��E�y`9���_jE�wj���8 �!�
endstream
endobj
62 0 obj
<<
/Size 63
/Root 1 0 R
/Info 59 0 R
/ID [<D0DE5E7D89EADD4DA09B2C6049C6F9E1> <221E9B4AFA953798F1C50210952E9A16>]
/Type /XRef
/W [1 3 2]
/Filter /FlateDecode
/Index [0 63]
/Length 208
>>
stream
x�-ЫR�Q൐�� ���Y�@����X�OD�'�AH4�S�d́����͞���9� ��B~������`�����������i�˭��hC	qy#c2l��2�<�����\��V&dR��޷�i�!�~=)ʬ��<�9{{'�a�IM�˒,?Co+�J&#�m�����:��+d���z�"_�}n�W���+s=17U�
�P�
endstream
endobj
startxref
100373
%%EOF
